 
Justering av protokollet från föregående sammanträde Protokollet från gårdagens sammanträde har delats ut .
Finns det några synpunkter ?
Herr talman !
Jag ser i protokollen att två ledamöter i går talade om försenade flyg till Strasbourg i måndags .
Jag skulle vilja tillägga att flyget från Amsterdams Schipol-flygplats också var försenat och senare blev inställt .
Vi omdirigerades till Basel-Mulhouse-flygplatsen .
Man talade om för oss att en buss skulle möte oss där när vi kom fram .
I själva verket dröjde det 45 minuter efter vår ankomst innan en buss anlände till flygplatsen .
Till slut kom vi hit , i måndags klockan 20.30 , efter att några av oss hade varit på resande fot i mer än tolv timmar .
Denna slags service och svårigheter för att komma till Strasbourg på en måndag är någonting ganska hopplöst .
Om den franska regeringen insisterar på att vi skall fortsätta att sammanträda i Strasbourg , kan den åtminstone se till att det när flyg omdirigeras till Basel finns bussar som kommer i tid för att möta de omdirigerade passagerarna , annars är det ganska meningslöst för oss att försöka komma hit på måndagar för att delta i arbete av något slag .
Jag undrar om detta kan föras till protokollet ?
Herr talman !
Jag var bokad på samma flygplan , och skäms över att behöva säga att det i detta fall handlade om KLM , vårt nationella flygbolag , och jag hoppas att det kan bli bättre nästa gång , även i fråga om samarbetet med ett annat flygbolag .
( Protokollet justerades . )
Herr talman !
Jag vill bara påpeka något som rör dagens föredragningslista .
I måndags beslutade vi att rådets förklaring med anledning av Genèvekonventionens 50-årsjubiléum skall skjutas upp .
Jag vill bara klargöra att det i dag endast handlar om övriga punkter på föredragningslistan , inte om Genèvekonventionens 50-årsjubileum .
Den punkten har skjutits upp till nästa sammanträde i mars .
Av misstag är punkten fortfarande upptagen på dagens föredragningslista .
Ledamot Swoboda , jag kan bekräfta det ni just sagt .
Det rör sig om ett tryckfel .
Den text som delats ut är felaktig , för det har beslutats att diskussionen skall senareläggas .
Herr talman !
Jag vill bara säga att jag när jag kom hit i morse noterade att två personer rökte utanför salen .
Lukten är fruktansvärt motbjudande !
Kan ni vara vänlig att göra någonting åt det ?
Personligen tror jag inte att jag kan göra det , men ni har rätt : vi måste försöka hitta ett snabbt sätt att lära upp dem som inte respekterar de förbud som vi själva har beslutat om .
När det gäller de försenade flygplanen och de problem som detta har ställt till , så skulle man kunna bilda en liten förening - jag vet inte riktigt hur liten - för dem som har haft svårt att komma till Strasbourg i tid för denna sammanträdesperiod , med uppgift att analysera hur många och vilka problem som faktiskt uppkommit .
 
Samstämmigheten mellan unionens olika politikområden och utvecklingspolitiken Nästa punkt på föredragningslistan är uttalanden av rådet och kommissionen - Samstämmigheten mellan unionens olika politikområden och utvecklingspolitiken .
Herr talman !
Det är en stor glädje för mig att i dag kunna vända mig till er här i kammaren i egenskap av rådets ordförande .
Jag vet att Europaparlamentets roll den närmaste tiden när det gäller behovet av att förstärka utvecklingspolitiken på unionsnivå är av stor vikt .
Mitt uttalande i dag har att göra med utvecklingspolitikens samstämmighet inom Europeiska unionen .
Jag kommer givetvis att låta kommissionen komplettera en del av mina kommentarer .
Jag vill börja med att betona det behov som vi alla inom Europeiska unionen har när det gäller att förena den extraordinära utveckling och de framsteg vi fått erfara i våra livsvillkor , främst tack vare den under de senaste årtiondena allt starkare teknologiska impuls som gynnat stora delar av världens befolkning vad gäller välstånd och förbättrade livsvillkor , med det faktum att vi samtidigt kan se att skillnaderna mellan en del regioner och geopolitiska områden i världen har ökat , vilket sätter det internationella stabilitetssystemet på spel och hotar freden .
Detta gör att vi alla måste följa vårt samvete och på bästa möjliga sätt försöka anpassa vår politik till målet om ökad stabilitet och större jämvikt mellan olika områden på vår planet .
Detta innebär att vi måste omvärdera utvecklingspolitiken som svar på globaliseringen av de ekonomiska och finansiella marknaderna .
Man har kunnat konstatera stora skillnader i marknadernas funktionssätt , vilket givetvis innebär att viktiga ändringar behöver göras , något som i sin tur ger utvecklingspolitiken nya möjligheter .
Vi står därför på tröskeln till ett nytt paradigm vad gäller utvecklingspolitik som , vilket jag gärna betonar , kräver att våra åtgärder koncentreras på fyra grundläggande aspekter : För det första , ett mera samstämmigt agerande mellan alla internationella aktörer på givarnivå , vi måste verka för större samordning , samstämmighet och samband mellan det humanitära biståndet och utvecklingspolitiken , vi måste få ett starkare multilateralt system , och vi måste uppmärksamma skuld- och finansieringsproblematiken .
Det kommer emellertid också att ställas nya krav på de länder som i dag tar emot stöd .
De måste bekämpa korruptionen , de måste styras av en demokratiskt vald regering , det vill säga grundläggande principer för en utveckling av landets politiska system , samtidigt måste de uppmärksamma sin egen politik och bekämpa fattigdomen .
En annan aspekt av utvecklingspolitikens nya paradigm har sin upprinnelse i behovet av att ha en mera integrerad syn på utvecklingen , den skall inte bara betraktas som ett stöd för tillväxten , då bör man hellre värdesätta andra typer av politik inom områdena för ekonomi , handel och investering , givetvis , men den har också sin upprinnelse i behovet av en mera integrerad syn på utvecklingen vare sig det gäller den globala politiken eller politiken i de olika givarländerna .
En tredje aspekt som jag skulle vilja betona när det gäller det nya paradigmet baseras på en målinriktad politik .
Sedan 1995 , efter att de främsta givarländerna på internationell nivå försökt komma överens om några viktiga uttalanden som gjordes i OECD : s kommitté för utvecklingsstöd , har man kunnat fastställa några viktiga mål för att leda och verkställa utvecklingspolitiken , må vara på nationell eller på internationell nivå .
Med dessa mål inriktar man sig på att halvera fattigdomen fram till år 2015 , må vara , som alla vet , genom att höja den obligatoriska skolgången eller kraftig sänka barndödligheten eller ingripa i den sociala välfärden så att man effektivt kan nå målet .
Detta skulle innebära att man tog bort den extrema fattigdomen för mer än en tredjedel av världsbefolkningen , vilket måste betraktas som något alldeles extraordinärt , men skall målet nås krävs säkerligen ett stort deltagande och ett kraftigt ingripande av hela det internationella samfundet Det här var den fjärde aspekten på den nya utvecklingsparadigm jag ville belysa : dagens utvecklingspolitik , särskilt de senaste årens utvecklingspolitik , styrs alltmer av globala frågor men det saknas ett starkt internationellt ledarskap .
De åtgärder som vidtagits av Förenta nationernas institutioner har starkt bidragit till detta , men så har även " Bretton Woods " systemet .
Det är värt att notera de mycket betydelsefulla impulser som Världsbanken har gett genom sitt dokument Comprehensive Framework och genom Internationella valutafonden .
Det är första gången en institution av det här slaget tar upp problemet om hur fattigdom skall avhjälpas som en central politisk fråga och öppnar en förbindelse , som fram till dess var otänkbar för en sådan institution , mellan skuldkvittning och fattigdom .
Det portugisiska ordförandeskapet har betonat att Europeiska unionen har ett stort behov av att förena sin mycket viktiga roll som huvudgivare på det internationella planet med en ledande och mera aktiv roll för att förnya utvecklingspolitiken på internationell nivå och åstadkomma bättre samordning mellan Förenta nationernas system och " Bretton Woods " systemet .
För att de skall vara möjligt att bearbeta Europeiska unionens roll i den internationella utvecklingspolitiken menar vi att vi först och främst måste vidta tre åtgärder .
För det första måste vi effektivisera utvecklingspolitiken .
År 1995 utvärderades som ni alla vet utvecklingspolitiken globalt och under det tyska ordförandeskapet kunde man lägga fram slutsatserna av denna globala utvärdering .
I de huvudsakliga slutsatserna betonar man vikten av en mera sammanhängande politik och ett allmänt strategiskt sätt att se på utvecklingsproblemen från Europeiska unionens sida .
Man betonar behovet av större samordning och kompletteringsmöjligheter mellan de olika politikområdena , och man måste också harmonisera och förenkla de organisationsformer som man i dag använder för att verkställa unionens samarbetspolitik .
Det finns också ett behov av att effektivisera hanteringen av stödet och på nytt gå igenom interventionsmekanismerna , och även utvärderingssystemet måste förstärkas och större öppenhet i förfarandet efterlyses .
En annan aspekt som är värd att belysa är behovet av kompletteringsmöjligheter mellan Europeiska unionen och medlemsstaternas politik .
Vi vet att en stor del av dagens stöd är ett resultat av medlemsstaternas nationella politik , stöd som inte alltid är kompletterande eller samordnade .
En stor del av den förspillan och ineffektivitet som Europeiska unionens stöd får vidkännas beror just på denna oförmåga att samordna och komplettera vad varje medlemsstat gör och vad Europeiska unionens institutioner föresätter sig att göra .
Vi menar att det är absolut nödvändigt att vi alla inom kort kan förstärka kompletterings- och samordningsmekanismerna mellan medlemsstaternas politik och Europeiska unionens politik .
Den tredje aspekten som är värd att belysa är en starkare och mera samstämmig politik , det centrala temat i dagens föreslagna debatt .
För det första så vet vi alla att det inte räcker med att förbättra villkoren för stödet och vi vet också att Europeiska unionen måste förbättra sina andra politikområden , så att utvecklingsmålen inte bara kan nås genom stödåtgärder och annan hjälp , utan först och främst genom att ha en mera integrerad syn på de politikområden som bidrar till utvecklingsmålen .
Som ni vet godkände rådet i juni 1997 en resolution , kommissionen lovade en utvärderingsrapport och det första betänkandet överlämnades till rådet i maj 1999 .
Redan här tas vissa samordningsaspekter upp , nämligen inom områdena för fred , livsmedel , fiske och migration .
Men vi väntar också på ett meddelande från kommissionen om samstämmighet tillsammans med ett meddelande om " Utvecklingspolitik " .
Den här debatten kommer givetvis under de närmaste månaderna , fortfarande under portugisiskt ordförandeskap , att berikas av det som kommissionen inom kort presenterar .
Samstämmigheten mellan olika politikområden kommer givetvis alltid att vara begränsad och en och annan motsats mellan dem är bara naturligt och utgör till och med en slags jämvikt och eftertanke mellan motsatta och konfliktskapande intressen , vilket ger liv och rörelse åt unionen , och att det bara är på det här sättet som det är möjligt att reglera motsatserna mellan de olika områdena .
Oberoende av detta vill vi understryka att bättre samstämmighet mellan olika politikområden inom Europeiska unionen , i nuläget och med den konjunktur vi har i unionen , innebär att vi noggrant måste överväga en del aspekter som har att göra med Europeiska unionens inre dynamik .
Vi vet att Europeiska unionen har en egen dynamik , i första hand baserad på Amsterdamfördraget , som förstärker den politiska dimensionen , något som tvivelsutan starkt berör budgeten för samstämmighet mellan politikområden och utvecklingspolitiken .
Vi måste också invänta regeringskonferensens arbete , se vilken väg man väljer för utvidgningen och hur långt Europeiska unionens inre dynamik inriktas på att förbättra samstämmigheten mellan politikområdena , främst utvecklingspolitiken , och om man också är beredd att inrätta lämpliga institutioner för ett sådant ändamål .
En annan aspekt vi måste begrunda när det gäller samstämmighet mellan politikområden är utvecklingspolitiken inom ramen för unionens utrikespolitik .
Vi vet att unionen ser på utrikespolitiken med andra ögon , vi vet att vi med inrättandet av Höge representanten , den snabba insatsstyrkan och centrumet för militär krishantering , har en hel del påtagliga bevis som vi inte får underskatta när vi tar itu med utvecklingspolitiken .
Det finns också aspekter som har att göra med den politiska dialogen , godkännandet av gemensamma ståndpunkter eller åtgärder , förberedandet av gemensamma strategier , den förebyggande diplomatin , utvecklingen av den regionala förmågan att förebygga och hantera krissituationer .
Alla de här aspekterna kommer givetvis när de införlivas och utvecklas att bidra till en bättre utvecklingspolitik inom ramen för Europeiska unionens utrikespolitik .
Vi kan säga att även på den här nivån , på Europeiska unionens nivå , måste utvecklingspolitiken inom ramen för utrikespolitiken gå samma väg som utvecklingspolitiken i många medlemsländer gjorde , det vill säga inom ramen för respektive lands utrikespolitik .
Ett sådant påstående förutsätter givetvis att man måste förbättra beslutsmekanismerna och de institutionella strukturerna med hjälp av GUSP , så att samordningen mellan de utvecklingspolitiska och utrikespolitiska instrumenten blir bättre .
I det här sammanhanget är vi övertygade om att vi måste lämna ett postkolonialt paradigm och övergå till ett genuint europeiskt paradigm för utvecklingspolitiken , eftersom vi vet att utvecklingspolitiken i ett europeiskt perspektiv har varit mycket beroende av en del länders politik och deras förhållande till den postkoloniala politiken .
En tredje aspekt att beakta är Europeiska unionens politik och medlemsstaternas politik .
Samstämmigheten mellan politiken på Europeiska unionens nivå förutsätter givetvis en bättre samordning av medlemsländernas politik och Europeiska unionens politik när det gäller utvecklingspolitiken .
Är det omöjligt att uppnå bättre samstämmighet mellan de nationella politikområdena så kommer det säkerligen att vara än svårare att tänka sig samstämmighet för Europeiska unionens utvecklingspolitik .
En fjärde och sista aspekt jag skulle vilja att ledamöterna begrundade när det gäller utvecklingspolitiken är rollen för rådet ( utvecklingssamarbete ) .
De senaste månaderna har man särskilt diskuterat dess roll i unionspolitiken .
Skillnaden mellan utvecklingspolitiken och annan politik på unionsnivå när det gäller förordningar är som vi alla vet flagrant - det räcker med att se hur svårt det var med EUF : s budgetering eller icke budgetering - och det är svårt att tro att vi kan få bättre samstämmighet mellan Europeiska unionens olika politikområden utan en mera aktiv och intervenerande roll från rådets ( utvecklingssamarbete ) sida när det gäller att bistå politiska beslut som uppenbart borde hanteras vid andra utvecklingsforum men som nu bearbetas av andra råd , av andra beslutscentrum , allt från Agrifin-rådet och rådet ( fiske ) till rådet ( miljö ) , och där rådet ( utvecklingssamarbete ) fram till nu inte har haft någon möjlighet att göra sin röst hörd eller på annat sätt ingripa .
Om rådet ( utvecklingssamarbete ) inte får spela en mera aktiv roll i den globala samordningen av politiska beslut , vilket direkt berör Europeiska unionens utvecklingspolitik som utformas vid sidan av olika beslutscentrum , kommer det säkerligen att bli mycket svårt att utveckla en mera samstämmig politik inom Europeiska unionen när det gäller utvecklingsmålen .
Vi välkomnar Europaparlamentets åsikter som säkerligen kommer att vara lämpliga .
( Applåder ) .
( EN ) Tillåt mig att först säga några ord om de framgångsrikt avslutade förhandlingarna mellan EU och AVS-länderna .
Jag skulle vilja påpeka att det var en mycket positiv upplevelse att delta i dessa förhandlingar .
Jag såg medlemsstater arbeta som ett lag , vilket verkligen var en underbar upplevelse .
Båda sidor var också mycket nöjda när det var över , inte bara för att det var över , utan för att vi alla visste att vi hade uträttat någonting tillsammans , EU och de 71 AVS-länderna .
Det är någonting som världen behöver , och det är en mycket bra signal inom ramen för hela globaliseringsdiskussionen .
Jag skall ange huvuddragen i några av de större nyheterna i det nya avtalet .
Vi tar uttryckligen itu med korruptionen ; vi upprättar en ram för att angripa problemet med invandring för första gången någonsin .
Vi främjar deltagarinriktade tillvägagångssätt , vi säkerställer att det sker samråd med det civila samhället om de reformer och strategier som skall stödjas av EU .
Vi riktar om utvecklingspolitiken till strategier för att minska fattigdomen .
Vi grundar fördelningen av biståndet inte bara på en uppskattning av varje lands behov , utan även på en uppskattning av resultaten av tidigare strategier .
Vi skapar ett investeringsorgan för att stödja utvecklingen i den privata sektorn .
Vi rationaliserar instrument och inför ett nytt system med rullande planering , vilket tillåter gemenskapen och mottagarländerna att regelbundet anpassa sina samarbetsprogram .
Vi decentraliserar det administrativa och , i vissa fall , det finansiella ansvaret till lokal nivå , med målet att effektivisera samarbetet .
Vi förbättrar den strategiska ramen för utveckling av handel och investeringar .
Vi ökar samarbetet på alla områden som är av betydelse för handeln , och här inbegrips nya frågor som arbetsnormer och kopplingen mellan miljö och handel .
Jag är säker på att ni efter Seattle kommer att uppskatta betydelsen av dessa avtal .
Tillåt mig att gå över till några av de viktigare punkterna .
För det första , avtalet om politiska frågor .
Det nya avtalet kommer att innebära att båda sidor förbinder sig att erkänna god skötsel av den offentliga verksamheten som en grundläggande och uttrycklig beståndsdel i partnerskapet , ett föremål för regelbunden dialog på ett område som åtnjuter gemenskapens aktiva stöd .
För det andra har ett nytt förfarande utarbetats för fall då kränkningar av de mänskliga rättigheterna , de demokratiska principerna och rättsstatsprincipen äger rum .
Jämfört med det nuvarande förfarandet , betonas de berörda staternas ansvar i större utsträckning enligt det nya förfarandet , och det tillåter större flexibilitet i samrådsprocessen , i syfte att få till stånd en effektiv dialog som leder till att åtgärder vidtas för att rätta till situationen .
I särskilt brådskande fall , då särskilt allvarliga kränkningar av någon av dessa oundgängliga beståndsdelar har ägt rum , kommer åtgärder omedelbart att vidtas , och den andra parten kommer att underrättas .
För det tredje har EU och AVS även enats om ett nytt speciellt förfarande som skall tillgripas vid allvarliga fall av korruption .
Detta är en verklig nyhet , både i EU-AVS-sammanhanget och då det rör sig om internationella förbindelser i allmänhet .
Detta förfarande kommer inte bara att tillämpas i fall av korruption där pengar från Europeiska utvecklingsfonden ( EUF ) är inblandade , utan också mer allmänt i varje land där EG är ekonomiskt inblandat och där korruption utgör ett hinder för utvecklingen .
Det är följaktligen inte begränsat till EG-verksamheter .
Detta är en mycket viktig aspekt , om man beaktar de offentliga finansernas kapitaliseringsförmåga .
Genom att ta med en sådan bestämmelse i partnerskapsavtalet , sänder EU och AVS-staterna tillsammans en tydlig och positiv signal , som utan tvekan kommer att uppskattas av europeiska skattebetalare och förhoppningsvis också av europeiska investerare .
Ett annat nytt ämne i AVS-EU-avtalet gäller in- och utvandring .
Vi har nått en balanserad överenskommelse om samarbete på detta område .
Denna nya dimension i partnerskapsavtalet speglar de riktlinjer som EU , i enlighet med Amsterdamfördraget och slutsatserna från Europeiska rådets möte i Tammerfors i Finland i oktober 1999 , har anslutit sig till .
Europeiska unionen åtar sig att utveckla och tillämpa en invandrings- och asylpolitik som grundar sig på principen om partnerskap med ursprungsländerna eller ursprungsregionerna .
Avtalet som har slutits med AVS-länderna bereder vägen för nya initiativ , särskilt om rättigheterna för tredje lands medborgare inom EU , och för åtgärder som underlättar deras integrering .
Vi enades även om bestämmelser för att ta itu med frågor som hör samman med illegal invandring .
EU och AVS-staterna kommer att inleda den process som har som slutmål att definiera , inom en ram som skall framförhandlas med vart och ett av AVS-länderna , sätten och medlen för att avvisa invandrare som uppehåller sig illegalt på någon av parternas territorium .
Här omfattas även personer från tredje land och statslösa personer .
Dessa mycket nydanande strategier erbjuder ett bra tillfälle att förbättra skötseln av den offentliga verksamheten .
Avtalet tillhandahåller också en bra ram för att stödja de ömsesidigt förstärkande effekterna av handelssamarbete och utvecklingsbistånd .
Vi har enats om en process för att upprätta nya handelsuppgörelser med vilka man eftersträvar att liberalisera handeln mellan parterna och för att formulera bestämmelser om handelsrelaterade frågor .
Vad beträffar tidsramen för handelsförhandlingarna , har vi tillmötesgått AVS-staternas önskemål .
Förhandlingar kommer att inledas senast 2002 .
Denna tvååriga förberedelseperiod kommer att användas till att stärka regionala integreringsprocesser och AVS-ländernas förmåga att genomföra handelsförhandlingar .
En sexårsperiod är planerad för dessa förhandlingar .
Vi kommer att ta hänsyn till AVS-ländernas ekonomiska och sociala begränsningar på två sätt : för det första genom att låta de ekonomiska reformerna och handelsreformerna åtföljas av strategier för mänsklig och social utveckling samt , för det andra , genom att hjälpa AVS-staterna att bli aktiva aktörer i det internationella ekonomiska handels- och ekonomisystemet genom kapacitetsbyggnad och samarbete i multilaterala forum .
Detta tillvägagångssätt kommer att leda oss till ett system som är fullt förenligt med WTO-systemet .
Ekonomiska aktörer kommer att vara mer benägna att upprätta närmare förbindelser med sina AVS-partner .
De inhemska och utländska investeringarna kommer att öka , och mer kunnande och teknik kommer att överföras , och allt detta kommer att stärka AVS-ländernas konkurrenskraft och underlätta deras gradvisa integrering i världsekonomin .
Dessutom kommer avtalen med EU att fungera som ett ankare .
De kommer att befästa de ekonomiska reformerna , på samma sätt som de nationella och ekonomiska reformerna kommer att stabiliseras av båda parters åtaganden enligt avtalen .
Den logiska grunden bakom detta nya tillvägagångssätt är också baserad på idén att en politik för öppen handel i samverkan med en politik för social utveckling kommer att leda till ekonomisk tillväxt och minskad fattigdom .
En annan viktig aspekt är förbättringen av EU : s handelsystem gentemot alla de minst utvecklade länderna , av vilka 39 faktiskt ingår i AVS-gruppen .
Denna process kommer att äga rum under de kommande fem åren och leda till att exportörerna i de minst utvecklade länderna år 2005 kommer att ha fritt tillträde till EU-marknaden för i stort sett alla sina produkter .
Vad beträffar storleken på nästa EUF , har EU lämnat sitt budgetförslag .
Det är baserat på principen om att förena behovet av att bibehålla en betydande summa finansiella resurser i en tid av begränsade officiella budgetar för utvecklingshjälp med behovet av att göra gemenskapens bistånd effektivare .
I dag är omkring 9,5 miljarder euro av tidigare EUF-medel oanvända .
EU har förbundit sig att engagera dessa återstående balanser , plus de nya EUF-medlen möjligt för gemenskapen att avsevärt öka de årliga flödet av åtagande- och betalningsbemyndiganden under perioden .
Vi går de kommande åren följaktligen inte in i en period med minskad aktivitet , vi går in i en period med ökad aktivitet .
Ett sådant åtagande nödvändiggör en djupgående reform av förfaranden och tillämpningsstrategier hos båda sidor .
Det finns en mycket påtaglig länk mellan reformprocessen i kommissionen i sig och vår förmåga att leverera på platsen , vilket är grunden för uppgörelsen med AVS-länderna .
Om vi går över till vår utvecklingspolitik , skulle jag vilja säga att det globala sammanhanget har förändrats drastiskt .
Marginaliseringen av många ekonomier , ökad fattigdom i världen , behovet av bättre hantering av det ömsesidiga miljöberoendet , flyktingströmmarnas destabiliserande effekter samt de oroande konsekvenserna av väpnade konflikter och pandemiska sjukdomar utgör alla stora bekymmer .
Det är inom denna föränderliga globala ram som vi måste placera oss själva .
Lyckligtvis får vi genom utvärderingar av EG-biståndet ett meningsfullt verktyg för att förbättra vår verksamhet och förhoppningsvis även anta de utmaningar som jag nyss har nämnt .
Om vi skall koncentrera oss på resultaten från utvärderingarna , skulle jag vilja nämna följande problem : målen i gemenskapens politik är för många och för vaga , vilket påverkar samstämmigheten negativt .
Detta beror på komplexiteten i våra egna strukturer , men även på de mycket påtagliga inkonsekvenserna mellan den sektorinriktade politiken och intressena i medlemsstaterna .
Kommissionen har ett biståndssystem som är för komplext och fragmentariskt vad beträffar instrument , förfaranden och institutionella mekanismer .
Politiken fastställs ofta mer på grundval av de instrument som finns tillgängliga än på grundval av strategiska mål och tydligt definierade prioriteringar .
Vi har för litet personal i förhållande till den biståndsvolym som vi förväntas förvalta .
I genomsnitt finns det i kommissionen 2,9 personer för att förvalta 10 miljoner amerikanska dollar i bistånd , jämfört med 4,3 personer i Världsbanken och mellan 4 och 9 personer i större medlemsstater .
Detta är ett verkligt problem : det finns för många finansiella instrument , vart och ett med sina speciella särdrag , och i synnerhet en rad olika budgetrubriker .
Detta är svårt att förena med behovet av ett effektivt förvaltningssystem .
För att bemöta och lösa dessa problem , måste gemenskapen inleda en effektiv dialog med medlemsstaterna och parlamentet .
Det är absolut nödvändigt att vi tar itu med frågan om samstämmighet på ett realistiskt och pragmatiskt sätt , vilket betyder att debatten måste föras inom den lämpliga institutionella ramen , det vill säga i rådet och i parlamentet .
Vi måste också göra någonting åt bristen på samordnade åtgärder bland de 15 medlemsstaterna själva , liksom mellan dem och gemenskapen .
Genom att koncentrera gemenskapens utvecklingspolitik på internationellt överenskomna mål och strategier , kommer vi att göra det lättare för oss att bättre komplettera medlemsstaterna .
Detta är i mångt och mycket också den linje som presenterades av minister Amado .
När vi talar om politik nu för tiden , inlåter vi oss i en konvergeringsprocess .
Detta är en del av lösningen .
Vi är i färd med att utarbeta nya riktlinjer för vår politik , och det är nödvändigt att vi identifierar prioriteringsområden för gemenskapens handlande .
Allt har blivit mer och mer komplext .
Det gäller även för utvecklingssamarbetet .
Ingen enskild givare har möjlighet att angripa hela spektrumet av frågor , vilket sträcker sig från makroekonomiska frågor till lagstiftningsramen eller från sektorinriktad politik till en mångfald nya gränsöverskridande frågor , som kön , miljö , god skötsel av den offentliga verksamheten samt institutionella reformer .
Det är viktigt att vi finner flexibla mekanismer som tillåter en uppdelning av arbetet i enlighet med de olika givarnas kunnande och kapacitet i varje utvecklingsland .
Detta bör ske på medlemsstatsnivå och leda till att en sektorinriktad politik för gemenskapens agerande utformas .
Det är dit vi vill komma .
För att identifiera EG : s prioriterade stödområden , måste man räkna med gemenskapens speciella särdrag i förhållande till medlemsstaterna och de internationella institutionerna .
Jag skall bara nämna några få av dessa : vår förmåga att förena utvecklingspolitik och handelspolitik samt att säkerställa samverkan mellan bistånd och ekonomiskt samarbete ; vår neutralitet och vårt försvar av övergripande gemenskapsintressen ; det faktum att vi utgör en " kritisk massa " och kan genomföra relativt stora projekt , jämfört med vad enskilda medlemsstater normalt kan genomföra .
Dessutom , vår närvaro på platsen : i grund och botten ser jag som vår största fördel själva det faktum att vi genom att vara ett framgångsrik regionalt samarbetsprojekt själva ses som en neutral , välkommen partner för detta experiment över hela världen - något som vi är ensamma om .
Det är nödvändigt att göra gemenskapens politik effektivare och att utveckla en mer funktionsduglig strategisk ram .
Det är denna dubbla utmaning som kommissionen måste anta , genom att under de kommande månaderna utarbeta ett förslag till ett uttalande om den övergripande politiken .
Vi kommer att starta en bred och öppen samrådsprocess för att höra alla de olika berörda parternas åsikter .
I mina ögon är denna process inte riktigt men nästan lika viktig som innehållet , och vi kommer att lägga ned alla våra resurser på att delta aktivt , och vi inbjuder alla till att delta .
Parallellt med detta har vi även satt igång med processen för att öka samstämmigheten och klargöra och föra upp till ytan , ut i offentligheten , de verkliga eller inbillade problem som finns i detta avseende .
Detta kommer att vara en pågående process , som jag ser som ett slags försök till en oavbruten kvalitetskontroll , och jag inbjuder parlamentet till att delta i detta fortgående försök för att förbättra samstämmigheten i vårt verksamhet .
Herr talman !
Först och främst vill jag tacka Amado för hans ord och även ett tack till Nielson .
Jag gläder mig också över att Amado talade om EUF .
Problemet ligger dock inte här , hos parlamentet , och inte heller hos kommissionen ; rådet måste ta steget att budgetera EUF , så egentligen borde den predikan hållas i rådet .
Herr talman !
Ett tack också till herr Nielson .
Han talade utförligt om det nya Loméavtalet , men det är dock inte det egentliga ämnet för förmiddagens sammanträde .
Vi ville tala om samstämmighet .
Det är ämnet .
Ända sedan början av 1990-talet har Europaparlamentet , Europeiska kommissionen och Europeiska rådet erkänt att det inte står så bra till med samstämmigheten i den europeiska politiken , i synnerhet på området utvecklingssamarbete och på andra politiska delområden i unionen .
Dessa problem har uppmärksammats ett par gånger tidigare , år 1992 , år 1995 och år 1997 .
Alla exempel finns i en resolution som ligger framför oss .
Själv har jag i många år ställt frågor om denna problematik .
1997 upptogs till och med politisk samstämmighet som obligatorisk i Amsterdamfördraget .
År 1998 avtalades dessutom att Europeiska kommissionen årligen skulle ge ut en rapport där det skulle anges vilka förbättringar som uppnåtts .
Men vad har vi sett sedan dess ?
Vackra ord , även så i dag , men ingen rapport .
Det är egentligen så galet att man inte kan tala om det .
Man erkänner att det förekommer motstridig politik .
Man formulerar gång på gång goda föresatser , men i själva verket händer ingenting .
Det är således riktigt att vi tar upp detta här i dag .
För att illustrera dessa motstridigheter vill jag ge ett par exempel .
Ett antal utvecklingsländer odlar sockerrör för sockerproduktionen .
Inom unionen produceras också socker , via sockerbetor .
För att förhindra att detta billiga socker från utvecklingsländerna konkurrerar med det dyrare sockret från EU sätter man en rejäl importavgift på detta rörsocker .
Konsekvensen är att exporten av rörsocker från de berörda länderna till unionen avsevärt begränsas .
Samtidigt ger vi oerhört mycket utvecklingshjälp till dessa länder .
En minister från en av de karibiska öarna som odlar sockerrör sade en gång till mig : Om ni helt enkelt släppte in vårt socker i Europeiska unionen , då skulle vi över huvud taget inte behöva er utvecklingshjälp .
Ytterligare ett sådant exempel : kakaon .
Europeiska unionen vill tillåta en andel på 5 procent för alternativa fetter i choklad för att harmonisera den inre marknaden .
Det skulle också kunna vara noll procent , vilket också skulle harmonisera den inre marknaden .
Om man sätter andelen till 5 procent , då kan man vara nästan säker på att det missgynnar hundratusentals små kakaoodlare i utvecklingsländer .
Ändå förefaller det gå i den riktningen .
Vad är det då egentligen som vi håller på med ?
Det är också ett typexempel på den politik som får våra medborgare att säga : vad håller Bryssel på med egentligen ?
Det förefaller som om det europeiska näringslivet är viktigare här än våra egna principer , vår egen samstämmighet och utvecklingsländernas intressen .
Det finns också chockerande exempel på området sanktioner och embargon .
Varför genomförs en oljebojkott mot Haiti och inte mot Burma , där en vald president sitter fängslad , ett parlament har skickats hem och en del av parlamentsledamöterna har satts i fängelse eller till och med har mördats ?
Varför genomförs ingen oljebojkott mot Sudan , där många strider äger rum , nota bene med vapen som betalas med pengar från de oljebolag som är verksamma i de områden där flyktingarna finns ?
Här handlar det helt klart om kolossala inkonsekvenser .
Vi har nu återigen fått höra ett vackert exempel av Nielson beträffande det nya Loméavtalet .
Om det nya Loméavtalet rätt och slätt träder i kraft utan att alla dessa inkonsekvenser tas bort från politiken , då bygger politiken på sand för att använda ett bibliskt uttryck .
Rådet har gång på gång gett exempel på var det inte står rätt till : inom jordbruket , inom handeln , inom konfliktförebyggandet , inom fredsoperationerna , inom fisket , inom migrationen , inom miljön .
Kommissionär Nielson !
Det vi sitter och väntar på är en bra rapport om dessa inkonsekvenser och ett antal konkreta förslag för att ta bort dessa inkonsekvenser från politiken .
Än en gång , annars kommer alla era vackra exempel , hela er vackra politik - och det säger jag också till statssekreteraren - att vara byggd på sand , och det kommer inte att bli mycket av detta .
Medborgarna tar upp detta med oss .
Vi har själva ända sedan 1992 sagt : detta är ämnet för denna debatt .
Jag hoppas att detta budskap går fram till er ordentligt , och jag hoppas verkligen att ni inom kort kommer med en rapport med åtgärder .
( Applåder ) Herr talman , ärade rådsordförande , ärade kommissionär , ärade kolleger !
Helt i min kollega Maij-Weggens anda tror jag att det finns ett stort antal företrädare här som alla verkligen vill ta upp detta ämne .
Vi talar om ett ämne som är av grundläggande betydelse för Europeiska unionen .
Låt mig börja med att mycket exakt ange vad det är vi debatterar här .
Artikel 178 , avdelning XX i det konsoliderade Fördraget om Europeiska unionen lyder som följer : " Gemenskapen skall beakta målen i artikel 177 då den genomför sådan politik som kan beröra utvecklingsländerna . "
Vilka är då de mål som all politik i Europeiska unionen skall beakta ?
I artikel 177 specificeras detta mål som " en varaktig ekonomisk och social utveckling i utvecklingsländerna , särskilt i de mest missgynnade bland dessa , en harmonisk och successiv integration av utvecklingsländerna i världsekonomin , kampen mot fattigdomen i utvecklingsländerna " .
Herr talman !
Detta är inte några mål utan förpliktelser , detta är artiklar , juridiska artiklar , som utgör en del av det rättsligt fastställda regelverket som de europeiska institutionerna och medlemsstaterna skall hålla sig till .
Varje artikel i regelverket får naturligtvis inte bara bedömas utifrån dess juridiska giltighet , utan också utifrån hur viktigt innehållet är .
Jag anser , och lyckligtvis många med mig , att principen om politisk samstämmighet är av största vikt för varje statsmakt som vill vara en trovärdig tjänare för sina medborgare .
Det är bara en trovärdig statsmakt som är pålitlig som kan tillvarata medborgarnas intressen .
Detta är viktigt för den tillit som samhället sätter till statsmakten , men också viktigt med tanke på ändamålsenligheten , för samstämmighet är ett krav för att våra begränsade medel skall kunna användas på ett effektivt sätt .
Vi får inte måla verkligheten mer rosenröd än den är .
Verkligheten är motsträvig .
Det är statsmaktens uppgift att hantera detta faktum med öppenhet och insyn , utan bakvägspolitik .
Statsmakten är förpliktigad att visa vilka dilemman den har och var , när och varför det finns problem med den politiska samstämmigheten i stället för att bara smussla undan allt detta .
Det är inte ett lyxproblem vi talar om här i dag : fattigdomsproblematiken i tredje världen är ett oändligt och ömmande problem som kräver seriös uppmärksamhet .
Naturligtvis bevakar vi från parlamentets sida våra medborgares intressen , men det ligger också i våra medborgares intresse att leva i en stabil internationell omgivning där man eftersträvar mänsklig värdighet .
Det är ett moraliskt intresse , ett säkerhetsintresse och i slutändan är det till och med av intresse för vår ekonomi .
Vem är det egentligen som vinner på att skattepengar från den europeiske medborgaren går till hjälp åt Namibia för att stödja den ekonomiska utvecklingen när de fattiga boskapsskötarnas ekonomiska driftighet i samma land samtidigt undermineras på ett dramatiskt sätt av stenhårda exportbidrag , betalade av samma skattebetalare ?
Vi låtsas som om det inte äger rum , men vi vet alla att det äger rum .
Ärade kolleger !
Det är inte vår uppgift som parlamentariker att sticka huvudet i sanden som en struts .
Den allmännyttiga politiska samstämmigheten är därför ett ansvar för kommissionen som helhet , för rådet och för Europaparlamentet .
Kommissionären för bistånd kan inte ta detta ansvar ensam , hur gärna vi än ser honom här och hör honom tala , vilket också gäller för rådet ( biståndsfrågor ) och parlamentets utskott för utveckling och samarbete .
Här behöver vi en övergripande taktik .
Efter den mycket klara och skarpsinniga redogörelsen av såväl Amado som Nielson på den punkten vill jag gärna tillkännage att vi verkligen ser fram emot kommissionens förslag om att göra politiken i sin helhet samstämmig .
Inte bara från kommissionär Nielson , utan från kommissionen i sin helhet .
Därför uppmanar vi kommissionen i denna skarpa och tydliga resolution att utveckla konkreta instrument .
Vi måste tydliggöra var det förekommer problem med samstämmigheten och göra en inventering för att se vad dessa problem består av .
Vi måste visa vilka problem vi löser och vilka vi ännu inte har löst .
Därför pläderar jag för ett samstämmighetsobservatorium som tydliggör detta .
Därför måste vi inrätta arbetsgrupper i kommissionen , i rådet , i parlamentet , som kan övervaka samstämmighetsprocessen .
Herr talman , mina damer och herrar kolleger !
Om taket hos våra grannar läcker kan vi ge dem grytor och pannor för att samla upp vattnet i , men naturligtvis är det mer ändamålsenligt att hjälpa till med att täta läckan i taket .
Fjolårets kris i kommissionen är i dag löst , men för närvarande bör kommissionen komma med en politik där vi får fullt stöd för en taktik , för en samstämmighet som parlamentet otvivelaktigt kommer att kräva i resolutionen inom kort .
Jag önskar kommissionären lycka till med sin kamp inom kommissionen och Amado lycka till inom rådet .
Herr talman , kära kolleger !
Låt oss säga det med en gång : när det gäller samarbetspolitiken är samstämmighet långtifrån en principfast sak .
Fördragen föreskriver att Europeiska unionen skall hjälpa utvecklingsländerna i deras utveckling , men det finns många snedvridningar av dessa förklaringar i fördraget , vilket andra kolleger har framhållit på ett mycket bra sätt .
Den första bristen på samstämmighet har att göra med att unionen och medlemsstaterna inte är samordnade i fråga om utvecklingspolitik .
Detta medför betydande funktionsbrister , eftersom vissa av gemenskapsprogrammen läggs ovanpå nationella program , i stället för att riktas till projekt som inte har fått någon uppföljning .
Vi får också komma ihåg att vissa medlemsstater i praktiken för en neokolonial politik , vilket inte på något sätt bidrar till utvecklingen i de länder som får en så kallad hjälp .
Den andra bristen på samstämmighet hänger samman med stödet till despotiska regimer .
Man förklarar att en god förvaltning och ett slut på korruptionen är ett obligatoriskt krav , men man fortsätter att ösa in hundratusentals euro på bankkonton i Schweiz , via ett antal statschefers plånböcker .
Den tredje bristen på samstämmighet är förknippad med de mänskliga rättigheterna .
Man säger sig vilja skydda dem .
Man uppmuntrar utvecklingsländerna att respektera dem .
Man röstar till och med igenom ett stort antal resolutioner för att fördöma varje kränkning av dessa rättigheter .
Man ansluter sig också till internationella protester och kampanjer .
Fast samtidigt låter man vapenhandeln utvecklas , utan att ens bry sig om att begränsa handeln med de mest avskyvärda vapen : till exempel truppminor .
Och man gör inte särskilt mycket för att verkligen förhindra kränkningar av de mänskliga rättigheterna .
Den fjärde bristen på samstämmighet i Europeiska unionens samarbetspolitik är följande : hur önskar ni bidra till utvecklingen genom att plundra naturresurserna hos dem ni hjälper ?
Det krävs att Europeiska unionen lämnar fisken till de lokala fiskarna , så att de kan försörja den lokala befolkningen , i stället för att vi systematiskt förstör havets resurser .
Vi måste överlåta råvarorna till lokala producenter , så att de kan förädla dem .
Och man skall bara inte tala om oljan , för vi känner tyvärr till vilken politik som grupper som Elf och Total bedriver i Afrika .
För att gå ännu längre , och detta blir kanske snart en femte brist på samstämmighet , kräver vi en respekt för den biologiska mångfalden , bland annat för att alla skall kunna producera med eget utsäde och för att bevara de naturliga rikedomarna .
Men samtidigt - och det fick vi se vid de senaste förhandlingarna - förpliktar man AVS-länderna att underteckna TRIPS-avtalen , trots att det finns en risk för att de utsträcks till att omfatta levande organismer .
En sådan utvidgning av avtalen skulle betyda döden för den biologiska mångfalden och en återgång till ett faktiskt slaveri för de småjordbrukare i Syd som utelämnas till de multinationella bolagen .
Däremot , och det är en sjätte brist på samstämmighet , försvarar man inte tillämpningen av de befintliga fördragen .
Å ena sidan röstar man igenom ett budgetanslag för aidsbekämpning , men å andra sidan gör man ingenting för att införa ett krav på obligatoriska licenser inom ramen för de nämnda TRIPS-avtalen , vilket trots allt skulle tillåta utvecklingsländerna att producera egna läkemedel och bromsa det blodbad som har orsakats av aids .
Vid förhandlingarna inom WTO fortsatte Europeiska unionen i samma anda - trots att Schwaigerbetänkandet redan i den andra punkten framhåller att den pågående avregleringen av handeln knappast gynnar de breda befolkningslagren i utvecklingsländerna , särskilt inte de allra fattigaste - genom att försvara avregleringen av handelsutbyten och avskaffa , om än med några övergångsår , de förmåner som har beviljats AVS-länderna , när vi egentligen borde ha stärkt detta system , särskilt för de allra fattigaste länderna .
Den åttonde bristen på samstämmighet är av ett politiskt och praktiskt slag .
Man säger alltid : tänk globalt , agera lokalt .
Ändå försummar man lokala utvecklingsaktörer genom att föredra att diskutera med de nationella regeringarna och subventionera de icke-statliga organisationerna i Nord , på bekostnad av lokala program och icke-statliga organisationer i Syd .
Jordbruket och miljön är exempel på ytterligare problem , där det också finns brister på samstämmighet som man skulle kunna peka på , för att inte glömma forskning , utvandring och hälsa .
Kort sagt , man påstår sig vilja hjälpa utvecklingsländerna men uppmuntrar ändå avregleringen av marknaderna , samtidigt som man medger att detta strider mot ett sådant mål .
Låt oss säga det än en gång : Europeiska unionens samarbets- och utvecklingspolitik är inte sammanhängande .
Å Verts-gruppens vägnar uppmanar jag således parlamentet , institutionerna och kommissionen att tillsammans försöka uppnå samstämmighet i vår politik .
Herr talman !
Jag uppskattar i allra högsta grad dagens debatt , inte bara för att utvecklingsfrågan rent generellt är viktig utan också för att den är så aktuell .
Seattle blev ett misslyckande och förbindelserna mellan nord och syd bevisar detta av flera skäl .
Sammanträdet i denna nordamerikanska stad visade klart och tydligt på stora olikheter och djupa orättvisor för världens fattigare länderna .
Just nu och givetvis influerad av detta misslyckande organiseras Förenta nationernas tionde konferens för handel och utveckling i Bangkok .
Under tiden slutfördes , som tidigare nämnts , de förhandlingar som kommer att avgöra Lomékonventionens framtid .
Det här räcker för att visa hur viktig den här frågan är .
Dessutom har vi nästa toppmöte , Europeiska unionen - Afrikanska enhetsorganisationen ( OAU ) , som man till sist kom överens om att hålla i Kairo i april .
Oavsett analys , även om den är ytlig , gör att vi tvingas dra den slutsatsen att något , eller mycket , håller på att gå snett med nord-syd relationerna , vilket också inkluderar Europeiska unionen och utvecklingsländerna .
Det räcker med att nämna att den kategori länder som kallas mindre utvecklade under de senaste 30 åren har ökat från 25 till 48 och utgör i dag 13 procent av mänskligheten .
De står dock inte för mer än 0,4 procent av exporten och 0,6 procent av importen i världen .
Man kan också nämna den olyckliga omständigheten att de rika ländernas statliga stöd till utvecklingsländerna har minskat med 23 procent sedan 1990 .
De nedskärningar som nyligen gjorts i gemenskapsbudgeten för detta räkenskapsår visar också på samma tendens , vilket ger en dålig och politiskt felaktig signal .
Den trovärdige Michel Camdessus , fortfarande direktör för Internationella valutafonden , bekräftade i det tal han höll i söndags att arbetet med FN : s handels- och utvecklingskonferens ( UNCTAD ) har inletts , och här vill jag citera att " det internationella samfundet ger med en hand och tar med den andra " .
Han syftade givetvis på utvecklingsländernas stöd till de mindre utvecklade länderna .
Vilken ironi att ett sådant uttalande kommer från den det kommer , men sanningen är att det var så han sade och att jag fick tillfälle att höra det .
Det stämmer väl överens med verkligheten och det föranleder mig att säga att vi måste tänka om och lansera nord-syd relationerna på nytt men i annan form .
Europeiska unionens roll måste förändras samtidigt som det är sant att främjandet av en ny och mera rättvis och jämlik världsordning varken kan eller får upphöra att vara ett strategiskt mål för unionen .
Därför måste vi reflektera över den globalisering som sker och se vilka mera grundläggande inriktningar och dominerande intressen som ligger bakom det hela och , särskilt i det här sammanhanget , beakta vilka skadliga konsekvenser detta får för de mindre utvecklade länderna .
Att ett nytt avtal slöts med AVS-länderna är ett faktum .
Det är i sig ett positivt faktum , särskilt om vi beaktar de påtryckningar som gjorts för att få ett slut på det hela och att många länder inte ville se en fortsättning .
Vi kommer tids nog att få möjlighet att mera djupgående analysera avtalets exakta lydelse .
Det är dock sant att de europeiska förhandlarna var blygsamma och inte nådde ända fram till det som vi så lägligt hade föreslagit , även om nu det nya avtalet innehåller nya och innovativa förändringar .
En bidragande orsak till detta har en del politiskt viktiga drag i det nya avtalet om intresseföreningar varit .
Avtalet är utan tvekan ett resultat av komplicerade förhandlingar där båda parter fick göra betydande eftergifter ; Europeiska unionen när det gäller god regering och handel .
Först och främst var det dock ett resultat av AVS-gruppens ansträngningar , som på ett påtagligt sätt fick ny drivkraft av Seattle .
Jag vill särskilt framhålla att det verkar som om vi börjar få ett nytt sätt att se på de här frågorna , främst när det gäller handel , något som var välbehövligt .
Avslutningsvis måste vi gå längre med vår politik för utvecklingsstöd till utvecklingsländerna .
När det gäller finans och budget , skuldbördan , stödet till känsliga sektorer som exempelvis livsmedel och humanitär hjälp eller utbildning och hälsa , men även inom områdena för miljö , investeringar eller tillgången på information och ny teknik , liksom inom handelssektorn .
Samtidigt måste vi garantera en fullständig samstämmighet mellan utvecklingspolitiken och andra politikområden inom gemenskapen , men även mellan den politik som varje medlemsland bedriver .
Vi får inte nöja oss med att fortsätta med något som i grunden har visat sig vara otillräckligt och felaktigt .
Herr talman !
Efter att ha lyssnat på rådet och kommissionen i dag , måste jag helt enkelt titta på min föredragningslista .
Jo , det står faktiskt " Samstämmigheten mellan unionens olika politikområden och utvecklingspolitiken " .
Vi har emellertid inte hört ett enda ord om det , vilket jag tycker är väldigt pinsamt .
Vi har väntat på en rapport om samstämmighet i åratal .
Den borde ha funnits här i skriftlig form i dag ; och efter att ha hört kommissionär Nielson tala , har jag inte så svårt att föreställa mig att han kämpar mot mycket starka , motstridiga krafter i kommissionen .
Jag vet att kommissionären själv har både starka och ytterst förnuftiga synpunkter om samstämmighet och jag hade gärna hört dem i dag .
Eftersom man i det gemensamma resolutionsförslaget föreslår en rad effektiva mekanismer för att säkra samstämmighet , vill jag under min mycket korta talartid inskränka mig till att nämna ytterligare en , nämligen att kommissionen också bör utvärdera ny , relevant lagstiftning i detta sammanhang .
I övrigt vill jag koncentrera mig på den katastrofala effekt som EU : s gemensamma jordbrukspolitik har på utvecklingsländerna .
Dumpning av nötkött i Sahel och Sydafrika , tomatpuré i Västafrika , mjölkpulver i Jamaica - exemplen är förhoppningsvis alla välkända .
De rammar åtminstone de berörda producenterna i AVS-länderna som måste förstöra sina produkter , eftersom de inte kan konkurrera med de statligt stödda produkterna från EU .
Europeiska skattebetalare bidrar med 40 miljarder euro om året till stöd för EU : s jordbruk .
Dessa pengar bidrar till att hämma utvecklingen inom jordbrukssektorn i utvecklingsländerna , som här utgör 69 procent av den totala arbetskraften mot 1,7 procent i EU .
Därutöver står jordbrukssektorn för 34 procent av utvecklingsländernas bruttonationalprodukt mot 5,3 procent i EU .
Här är det varken fråga om samstämmighet eller anständighet .
Varför vill varken rådet eller kommissionen erkänna det ?
Herr talman !
Hur man kommer fram till policybeslut är sannerligen av grundläggande betydelse .
Storbritanniens premiärminister och utrikesminister gjorde i går uttalanden om sin hållning i frågan om röstsystemet i rådet .
De påpekade att befolkningen i Förenade kungariket , Frankrike och Tyskland för närvarande med bred marginal överstiger befolkningen i de övriga länderna i Europeiska unionen .
De drog därefter slutsatsen att befolkningsstorleken bör avspeglas i röstsystemet och att Storbritannien inte kommer att ge upp sitt veto .
Diskuteras denna fråga i rådet ?
Är rådet berett att behålla ett demokratiskt veto som baseras på befolkningsstorlek , eller går det fortfarande i riktning mot ett röstsystem med enkel majoritet av rådsledamöterna , i stället för ett röstsystem som speglar den befolkning i Europa som de demokratiskt företräder ?
Har Förenade kungarikets företrädare gett uttryck för sitt beslut och förslag för rådet , och vilken , om någon , hänsyn har man tagit till det ?
Då denna röstsystemsfråga är livsviktig för unionens demokratiska framtid , bör det utan tvekan ges högsta prioritet .
Hur besluten fattas är av grundläggande betydelse .
Herr talman !
Jag tackar rådet och kommissionen för deras uttalanden denna förmiddag , men jag kommer att koncentrera mig på frågan om samstämmigheten mellan politikområden , eftersom det är vad föredragningslistan säger att vi skall tala om .
Trots att jag håller med om behovet av att hålla en debatt om samstämmigheten mellan unionens olika politikområden och utvecklingspolitiken , är jag inte säker på att det i dag är rätt tillfälle att hålla den .
Rådets uttalande gav mig emellertid hopp om framtiden .
Det är ganska uppenbart för mig , som en person som har specialiserat sig på utvecklingspolitiken , att det finns många områden där bristen på samstämmighet på ett dramatiskt sätt påverkar utvecklingsnationerna .
Jag skall strax ge några exempel .
Jag påminner emellertid kammaren om att man i juni 1997 i en rådsresolution erkände det faktum att det finns en allvarlig brist på samstämmighet mellan vissa av EU : s politikområden och dess utvecklings- och samarbetspolitik .
Detta följdes av en begäran från rådet till kommissionen om att tillhandahålla en årsrapport , och det var tänkt att den första av dessa skulle diskuteras 1998 .
Vi väntar fortfarande på den första rapporten , och det är därför jag anser att denna debatt hålls för tidigt , då kommissionen inte hade mycket att säga om samstämmighet denna förmiddag .
De områden som identifieras av rådet är specifika områden där det är särskilt viktigt med samstämmighet mellan olika politikområden , som till exempel fredsbyggande , konfliktförebyggande och konfliktlösning , livsmedelssäkerhet , fiskeripolitik samt invandring .
Några av dessa frågor har diskuterats grundligt .
Jag tycker personligen att frågor som fredsbyggande och konfliktförebyggande och konfliktlösning i mångt och mycket bör hanteras av de afrikanska statsöverhuvudena , med kapacitetsstöd från Europeiska unionen och Afrikanska enhetsorganisationen ( OAU ) i rollen som skiljedomare .
De frågor som verkligen berörs av bristen på samstämmighet återfinns på områden som jordbruk , handel , miljö och biologisk mångfald , men häri ligger det verkliga problemet : det rör sig om extremt känsliga politikområden , i Europeiska unionen i allmänhet och i detta parlament i synnerhet .
Ledamöterna i denna kammare skulle ha olika åsikter , även inom samma politiska partier , beroende på a ) vilket land de kommer ifrån eller b ) vilket utskott de sitter i .
Det finns områden mellan vilka jag , som ledamot av utskottet för utveckling och samarbete , skulle vilja se samstämmighet som förmodligen skulle förskräcka vissa av ledamöterna i utskottet för jordbruk och landsbygdens utveckling eller i fiskeriutskottet .
Som ett exempel på bristen på samstämmighet kan man anföra , vilket Sandbæk gjorde , exporten av mjölkprodukter till Jamaica till priser långt under produktionskostnaderna i landet , vilket nästan ödelade den jamaicanska mejeriindustrin .
Vi exporterar nötkött till södra Afrika , till Namibia och Sydafrika , som sedan säljer sitt inhemska nötkött till Swaziland , så att Swaziland kan fylla sin exportkvot tillbaka till Europeiska unionen .
Kom också ihåg att vissa länder blockerade ett handelsavtal med Sydafrika i fyra år .
Om vi bara importerar råmaterial från dessa utvecklingsländer , i stället för att tillåta dem det mervärde som det medför att färdigställa varorna i det egna landet , förvägrar vi dem just den fattigdomsbekämpning som vi har satt som vår huvudprincip då det gäller hjälp till utvecklingsnationerna .
Det förvånar mig inte att kommissionen har svårigheter att framställa ett grunddokument för en diskussion om en hållbar och social utveckling .
Det finns ett naturligt motstånd i tredje världen mot allt som skulle sänka levnadsstandarden och skapa ytterligare arbetslöshet .
Jag önskar kommissionen lycka till i sin ansträngning att framställa detta grunddokument .
Herr talman !
Den här förmiddagens debatt är en mycket viktig debatt .
Jag vill därför tacka kommissionen och rådet som har uttalat sig om samstämmigheten mellan unionens olika politikområden och utvecklingspolitiken , för det är ett bevis på att det finns en vilja att göra politiken effektivare i det avseendet .
Om vi inte gjorde något mer än att konstatera bristen på samstämmighet i vår politik skulle det skapa en stark frustration hos oss och det är enbart negativt .
På samma sätt som för styrkeförhållandena som studeras inom den elementära fysiken är det ingen mening med att införa politikområden som motverkar varandra .
Resultatet av ett sådant absurt spel är inte lika med noll , utan det skulle till och med skapa ett negativt värde , bestående av de materiella , finansiella och mänskliga resurser som har slösats bort på en värdelös satsning .
Ett negativt värde som inom politiken multipliceras med det antal resultat som inte kan uppnås varje gång en åtgärd häver de effekter som en annan åtgärd hade avsett att ge .
I dagens globaliserade värld är det en uppenbart faktum .
Det finns inte heller några gränser för gemenskapens politikområden .
Därför gläder det mig att kommissionen och rådet åter visar intresse för samstämmigheten mellan gemenskapens politikområden och att de , förutom de nationella politikområdenas kompletterande av varandra och gemenskapens politik och samordningen av kommissionens tjänster , har för avsikt att anpassa partnerskapspolitiken till utvecklingen inom Europeiska unionen .
Såväl kommissionen som rådets portugisiska ordförandeskap uttalar i sina arbetsplaner en önskan om samstämmighet mellan de politikområden som i stor utsträckning påverkar utvecklingsländerna , men utan att specificera vilka konkreta åtgärder denna samstämmighet skall ta sig uttryck i .
Båda institutionerna klargör vilka områden detta koncept främst bör tillämpas på .
Det framgår till exempel av kommissionens långsiktiga planering att målet i form av en hållbar utveckling bör ta sig uttryck i en stark solidaritet , med stöd av en handelspolitik som beaktar de gemensamma intressena .
Kommissionen hänvisar till ett mycket viktigt område , nämligen handelspolitiken .
Vi i parlamentet vill lägga till politikområden med stöd till utvecklingen , jordbruket , fisket , migrationen , unionens roll i de internationella finansinstituten , utrikespolitiken och säkerhetspolitiken och stödet till strukturanpassningen .
Rådet - det påpekade Luis Amado i morse - har redan vid flera tillfällen uttalat sig om behovet av samstämmighet - senast , och det stämmer , i november 1999 och även vid andra tillfällen , så som på rådsmötena för utveckling i maj 1999 och i juni 1997 - men utan några konkreta resultat .
Eftersom vi håller med om det han sade - som är av stor betydelse -är det inte mycket rådet för utveckling kan säga , precis som någon av föregående talare påpekade .
Däremot vill vi som parlament föreslå - och det framgår av resolutionen - att en arbetsgrupp för utbyte av tjänster tillsätts bestående av de ansvariga för alla nämnda politikområden , samt att ett observatorium inrättas för samstämmigheten mellan gemenskapens olika politikområden , där effekterna på varje område i utvecklingsländerna och länderna sinsemellan kan förutspås .
Vi vill i själva verket vara realistiska och vi är medvetna om att det för att vi skall uppnå målen med en samordning , en komplettering och det mest omfattande som vi nu håller på att behandla - samstämmigheten kommer att krävas en mer genomarbetad politik än den vi för närvarande har inom Europeiska unionen .
Låt oss hoppas - och det gör vi - att vi kommer att följa förändringens vindar från regeringskonferensen , från reformen av kommissionen - som även kommer att påverka utvecklingstjänsterna - , under denna nya mandatperiod med siktet inställt på en utvidgning för att skapa en mer samstämmig union .
Därför hoppas vi att kommissionen i den rapport som kommer att läggas fram inför parlamentet om den globala politiken även tar upp frågan om samstämmighet för en effektiv användning av gemenskapsresurserna och den konkreta förvaltningen av de offentliga intressena .
Herr talman !
Jag vill också gärna tacka rådet och kommissionen för deras redogörelser och i likhet med andra beklaga att samstämmighetspolitiken inte kommit mer i fokus .
Vi som sitter här i parlamentet tvivlar emellertid inte en sekund på vad som är orsaken till det .
Jag vill därför gärna ta upp något mer allmänt och inleda med ett par , tycker jag själv , beskrivande siffror .
I början av 1800-talet var realinkomsten per invånare i världens rikaste länder tre gånger högre än i de fattigaste länderna ; 1900 var den tio gånger högre och 2000 var den 60 gånger högre .
Det finns inga tecken på att denna utveckling kommer att vända ; tvärtom ser det ut som vi är inne i en exponentiell kurva som gör skillnaderna ännu större .
Det visar följande siffror : Inkomstklyftan mellan den rikaste och den fattigaste femtedelen var 1960 30 : 1 , 1990 60 : 1 och 1997 74 : 1 .
Dessa siffror härrör från perioden före Internetrevolutionens början .
Med andra ord : Det behövs enorma framsteg inom utvecklingspolitiken om inte de rika länderna , inklusive EU-länderna , skall bygga upp murar kring sig för att förhindra invandring i stor skala .
I den globala byn kommer de stora skillnaderna i världen inte längre att tolereras av den fattigaste delen av byn .
Vid en eller annan tidpunkt blir det uppror , och det är helt berättigat .
Jag vill därför uppmana rådets ordförandeskap att så snabbt som möjligt inleda den utlovade debatten och framför allt avsluta den , så att vi alla , inklusive Europas medborgare , kan förstå vad globaliseringen innebär och så att vi inser att ett centralt element blir genomgripande åtgärder på utvecklingsområdet vad gäller vårt utvecklingsbistånd och nivån på detta - vi ligger långt från de utlovade 0,7 procent som skall vara ett genomsnitt i EU .
Det kan vara så att andra är värre , men det hjälper inte oss .
Vi skall dock framför allt ge länderna möjlighet att handla med oss .
Såvitt jag hörde - men jag kan ha missat något - nämndes ordet handel över huvud taget inte i rådsordförandens tal .
Till kommissionären vill jag bara säga att jag hoppas det lyckas att få igenom hans förslag i kommissionen och medlemsstaterna , och jag vill också be kommissionären att ge några konkreta exempel på särintressen som inte bara blockerar i kommissionen , utan också i medlemsstaterna .
I övrigt vill jag gärna säga att jag tror att det mest effektiva skulle vara om parlamentet krävde att få ett förslag från både rådet ( utvecklingssamarbete ) och den kommissionär som är ansvarig för bistånd , så vi kanske fick en utgångspunkt för diskussioner istället för att kräva ett förslag från alla regeringarna och från hela kommissionen - det resulterar knappast i något positivt .
Jag skall avsluta med några ord om Internetrevolutionen .
Precis som kommissionär Liikanen reser runt och säger , så har vi ett försprång på mobilområdet här i Europa .
Låt oss utnyttja detta inte bara till förmån för de egna medborgarna , utan också till nytta för utvecklingsländerna .
Denna teknik möjliggör just de stora framsteg som behövs , och här kan EU bestämma dagordningen , prägla utvecklingen och leva upp till sitt globala ansvar .
Herr rådsordförande , kolleger , kommissionär Nielson !
Utan tankemässig samstämmighet på de olika områdena inom politiken går det inte , om man vill att utvecklingspolitik faktiskt skall leda till förbättringar .
Jag kan ju inte å ena sidan bygga upp något med ena handen för att strax därpå riva ner det igen med den andra !
Tyvärr måste man konstatera att en stor del av EU-politiken lider brist på just denna samstämmighet .
Detta gäller i alldeles särskild utsträckning jordbrukspolitiken .
För ännu i dag hindrar Europeiska unionen genom sin aggressiva exportpolitik och sin marknadsisolering utvecklingsländerna a ) i deras utveckling av ett självständigt jordbruk b ) att på ett skäligt sätt vara representerade med sina produkter på våra marknader .
Det är en jordbrukspolitik som ju inte bara skadar de små och medelstora producenterna i dessa länder , utan även tillverkarna i Europeiska unionen .
De spelas ut mot varandra .
Detta måste äntligen bli sagt och tas på allvar .
När jag ser , herr Armado , att det i ett land som Brasilien med en yta på över 8 miljoner km2 , som vid det här laget måste importera baslivsmedel , fortfarande finns nästan 40 miljoner undernärda och svältande människor , då måste jag säga att även detta i någon mån har att göra med hur vi driver vår jordbrukspolitik i och med att vi använder sojan därifrån för att producera våra nötköttsberg som vi i sin tur lägger på lager i kylhus !
Här ser vi tydligt att politiken måste förändras , men naturligtvis att det måste till förändringar till förmån för regionala strukturer även i utvecklingsländerna .
I framtiden kommer det vidare att vara avgörande vilken politik Europeiska unionen driver i Världshandelsorganisationen just till förmån för länderna i söder , på vilket sätt unionen vill ge dem en röst , ett rimligt medbestämmande där , och givetvis även i vilken mån Europeiska unionen öppnar sina marknader för dessa länder .
För inte kan det gå an att vi fordrar ett ömsesidigt öppnande av marknaderna i de här länderna , i just U-länderna , medan vi själva murar vidare här i Europeiska unionen .
Inte heller de handelsrelaterade regleringarna i TRIPS-avtalet ( Avtalet om handelsrelaterade aspekter på immateriella rättigheter ) går just dessa länders resurser till mötes .
För då måste de återigen betala dyrt för sina basprodukter här , som vi först tar patent på .
Låt mig ta upp ännu en punkt om samstämmigheten här i kammaren !
Ofta röstar man i de mest skilda utskott och även här i plenum , vilket inte direkt visar på samstämmighet , vilket inte överensstämmer med utvecklingspolitiken .
Därför borde utvecklingspolitiken vara ett tvärsnittsområde för alla utskott och inte som nu diskuteras bara en gång om året , just när det råkar vara opportunt .
Även politiken i de 15 EU-staterna måste samordnas på motsvarande sätt , för det går inte an att nationella intressen får fortsätta puttra med i den utvecklingspolitiska budgeten och att utvecklingsbiståndet kopplas till villkor som exempelvis : Köper du mina vapen så får du mer utvecklingsbistånd !
Så kan det inte få se ut i framtiden .
Mer samstämmighet är absolut nödvändig , det gäller inte bara Europeiska kommissionen och unionen , utan även oss här i kammaren !
Herr talman !
Rapporterna ger en redogörelse , men vittnar emellertid även om den växande inkonsekvensen i unionens och medlemsstaternas utvecklingspolitik .
När man konstaterar att bekämpandet av fattigdomen är den gemensamma nämnaren , då är detta snarare önskan än verklighet .
Faktum är att antalet fattiga människor de senaste 20 åren inte har minskat , utan ökat till 1,4 miljarder .
Ett ärligt bokslut för nord-syd-politiken kommer inte undan det faktum att glappet mellan de fattigaste och de rikaste länderna har vidgats än mer .
I stället för att beteckna detta som en direkt följd av den nyliberala politiken understryker man nödvändigheten av att tydligare definiera begreppet " god statlig skötsel " för utvecklingsbiståndet .
Jag undrar dock , med vilken moralisk rätt och med vilka anspråk skall detta göras när de fordrade kriterierna demokrati och rättsstatlighet kränks också i EU : s medlemsstater ?
Korruptionen blomstrar , svarta partikassor byggs upp , och EU-kapital leds förmodligen in i valkampskassor .
Att vi är kritiska mot oss själva är nu en förutsättning för att vi skall kunna fastslå reella kriterier .
Man skall heller inte glömma bort att unionens medlemsstater inte är i närheten av att avsätta 0,7 procent av bruttonationalprodukten till utvecklingsbistånd , tvärtom avlägsnar man sig alltmer från detta mål .
Vidare anser jag att det är beklagansvärt att det i rapporten inte spills ett ord på rustningsaffärer , andra kolleger har redan tagit upp detta .
Därmed gör industriländerna i förening med de härskande klasserna i flera AVS-länder inte bara våldsamma vinster , utan det sätts också igång ett fruktansvärt kretslopp som vi inte får glömma bort .
Först levereras vapen , sedan bryter det ut våldsamma konflikter , tills slutligen trupper från de vapenlevererande staterna sätts in , och så börjar allt om från början igen .
I Corries betänkande vill jag särskilt stödja konstaterandet att det finns anledning för oss att ge akt på rättvis behandling av Kubas medlemsansökan till AVS-länderna .
Där poängteras de förändringar som visar sig i inledningsskedet .
Vi bör inte följa USA , utan mer utgå från våra egna ställningstaganden och inte sätta upp nya , högre hinder .
Herr kommissionär , att kräva och skildra den politiska samstämmigheten är bra .
Men den vill även komma till uttryck i kommissionens politiska samverkan med parlamentet , och här tror jag att vi har stora uppgifter framför oss , som jag kommer att bidra till att utföra .
Herr talman !
" Det står illa till med Europeiska unionens utvecklings- och samarbetspolitik . "
Det är bara ett exempel på ett citat från en tidningsartikel förra veckan om unionens utvecklingspolitik .
Det är inga nya tongångar .
Även om vi i Europa försöker att göra något i fråga om utveckling och samarbete tvivlar man på dess effektivitet och kvalitet .
Förhoppningar om förbättring hotar att försvinna om kommissionen fortsätter att vägra se sig själv i spegeln .
Varför spreds inte den kritiska rapporten om sammanhanget i utvecklingspolitiken externt ?
En viktig slutsats i denna rapport avsåg den interna stridigheten om den europeiska politiken .
Det är i synnerhet på handels- och jordbruksområdet som den europeiska politiken står i strid mot utvecklingspolitiken .
Vi lyckas helt enkelt inte att ge ett seriöst bidrag till utvecklingen i de minst utvecklade länderna .
Allt detta har att göra med skillnaderna i synen på utveckling och samarbete mellan olika länder inom unionen .
Vi får inte längre betrakta utveckling och samarbete som instrument för externa och utrikes förbindelser , utan som självständigt politikområde .
Jag förespråkar en öppen , solidarisk och effektiv utvecklingspolitik .
Så länge en europeisk taktik i fråga om utvecklingspolitiken förorsakar mer ineffektivitet och mer slöseri med pengar är det tillrådligt att tilldela medlemsstaterna en stor roll .
Slutligen vill jag be kommissionen att skicka över det dokument som jag talade om så snabbt som möjligt , så att vi på ett konstruktivt sätt kan hjälpa till i tankearbetet med att hitta möjliga lösningar .
Herr talman , herr kommissionär , ärade kollegor !
Jag tycker att initiativet är lämpligt och meningsfullt .
Som mina kollegor redan har nämnt så står vi ofta inför mycket motsägelsefulla situationer där vi å ena sidan försöker föra fram utvecklings- och samarbetspolitiken och å andra sidan det som vi omintetgör genom annan sektoriell politik med motsatta intressen när det gäller samma länders utveckling .
Vi talar inte bara om den konkreta effekten av vår gemenskapspolitik , turism , miljö , jordbruk , fiske , industri .
Vi talar i mera allmänna ordalag , vilket är betydligt allvarligare , om motsättningar mellan vår ekonomiska och kommersiella politik och vår försvarspolitik .
Med andra ord , många motsägelsefulla situationer .
Jag menar att motsättningarna inom gemenskapspolitiken i själva verket inte är så allvarliga .
Då är det allvarligare det som sägs om vissa mål och industrier i en del medlemsländer .
Vi måste vara medvetna om detta .
Vi antar ofta resolutioner om fredsprocesser i andra delar av världen , som till exempel nyligen med Indonesien , vilket är himmelsskriande .
Efteråt kunde vi konstatera att det faktiskt fanns vissa länder i Europa som försåg dem med vapen och krigsmateriel .
Detta är för mig det mest motsägelsefulla i den här frågan , betydligt allvarligare än det motsägelsefulla i den sektoriella politikens oförenlighet , som också finns .
Visst vet vi att det finns motsättningar mellan varje lands politikområden .
Det är normalt .
Även på unionsnivå måste vi vara medvetna om att sådana motsättningar finns mellan olika gemensamma politikområden , i det här fallet utvecklingspolitiken .
Vi måste veta att motsättningarna finns och försöka minimera dem .
Målet att minimera motsättningarna är ett klokt och lämpligt mål och som presentationen av den här resolutionen grundar sig på .
Idén att inrätta en myndighet för att se hur denna samstämmighet utvecklas tycker jag är bra .
Verksamhetsområdet skall inte enbart begränsas till gemenskapspolitiken , utan det skall också omfatta politiska åtgärder vidtagna av medlemsländerna , inklusive ekonomiska gruppers aktioner , vilket jag tycker är viktigt .
Myndigheten skall årligen utarbeta en rapport om utvecklingen och effekterna av politiken i fråga och vad som därav kan härledas .
Den viktigaste frågan , enligt min mening , har jag lämnat till sist , en fråga som jag tror skall registreras och godkännas av parlamentet .
Vårt mål att minimera motsättningarna mellan utvecklings- och samarbetspolitiken och övriga politikområden måste vara ett giltigt mål inte bara inom Europeiska unionen utan också på internationell nivå tack vare den allt starkare globaliseringen av ekonomin .
Vill vi ha en rättvis världshandel måste den här principen tas med vid Världshandelsorganisationens nästa multilaterala förhandlingsrunda .
Det skulle nämligen vara motsägelsefullt om Europeiska unionen påförde sig själv en benhård princip , må vara rättvis , och att Förenta staterna eller annan stormakt sedan skulle göra det motsatta och utnyttja den .
Därför är det både rättvist och fundamentalt att den här principen klargörs vid Världshandelsorganisationens nästa runda .
Herr talman !
Generaldirektören för Generaldirektoratet för bistånd har sagt att det att framställa en rapport om samstämmigheten mellan EU : s politikområden och utvecklingspolitiken innan vårens dokument om själva utvecklingspolitiken läggs fram , är som att spänna kärran för hästen .
Det spelar ingen roll att kravet på kommissionen att framställa en årsrapport , ett krav som tydligt formulerades i rådets resolution , bara har resulterat i ett " icke-dokument " , det verkliga problemet här är att denna häst , samtidigt som fattigdom ökar i världen , stretar på uppåt medan kärran med EU : s andra politikområden är så tung att utvecklingspolitiken i själva verket sakta dras bakåt .
Gång på gång glöms utvecklingspolitiken bort , eller så kommer man att tänka på den i efterhand , när Europeiska unionens stora politikområden behandlas .
Ta det nya chokladdirektivet , som visar att EU-länderna spenderar mer på choklad varje år än på utvecklingsbistånd .
Det har inte gjorts någon lämplig bedömning av utvecklingsaspekterna i detta direktiv , som producentländerna , av vilka 90 procent är våra AVS-partner , uppskattar skulle kunna minska kakaoodlarnas inkomster med minst 15 procent .
Ta fiskeavtalen , där vi medger att den nuvarande fiskeripolitiken inom EU : s vatten är ohållbar .
Samtidigt förhandlar vi om samarbetsprojekt som skulle ge Europas storskaliga fiskefartyg ökat tillträde till utvecklingsländernas vatten , på bekostnad av arbetet för 190 miljoner personer som ägnar sig åt småskaligt fiske i dessa länder runt om i världen .
Ta handelsavtalen .
Som Nielson sade i förmiddags angående Lomé , gäller det prioriterade tillträdet enbart " i stort sett alla de minst utvecklade ländernas produkter " .
Med andra ord , när EU : s kommersiella intressen berörs , lägger man eventuella hänsynstaganden om fattigdom åt sidan .
Mot bakgrund av vår hållning i Seattle , varför råder det en sådan tystnad kring EU : s misslyckande att genomföra de handelsförmåner för utvecklingsländerna som redan har överenskommits inom ramen för GATT , inbegripet handelsförmåner för den viktiga textilsektorn ?
Vad gäller den gemensamma jordbrukspolitiken ( GJP ) , den största boven i dramat , har ingen bedömning gjorts av effekterna på utvecklingspolitiken av GJP-reformerna i Agenda 2000 .
Alla känner vid det här laget till skandalen med exportbidragssystemet , som ledde till att 54 000 ton nötköttsöverskott dumpades på västafrikanska marknader , vilket gjorde att priserna för de lokala boskapsuppfödarna halverades .
Det finns i dag ett nöttköttslager på 300 000 ton .
Vem står i tur att få benen undanslagna ?
Jag välkomnar Amadeus uttalande i förmiddags , i vilket han erkände svårigheterna med EDF-medlens icke-budgetisering , i vilket han uppmanade rådet ( utvecklingssamarbete ) till att spela en aktivare roll och i vilket han begärde att utvecklingsprioriteringarna skall bli centrala i EU : s framväxande gemensamma utrikes- och säkerhetspolitik .
Jag välkomnar även rådets förklaring från 1992 , dess resolution från 1997 och de successiva ändringarna i Fördraget om Europeiska unionen .
Åtgärder har bara inte vidtagits .
Det är därför vi vill ha årsrapporter , en årlig intern grupp för enheterna och ett klagomålsförfarande , för att säkerställa att åtgärder verkligen vidtas .
Jag ber herr Nielson att i sin sammanfattning direkt ta upp dessa punkter i resolutionen .
Herr talman !
Jag skulle vilja begränsa mig till förhållandet mellan utveckling och samarbete å ena sidan och jordbruk å andra sidan .
Under de senaste åren har en ansenlig del av fonderna gått till utveckling av jordbruk och boskapsskötsel , och då framför allt i Loméländerna .
Resultaten är inte direkt vad vi hade förväntat oss .
Vad skulle kunna vara orsaken till detta ?
Jag tror att orsaken i första hand måste sökas i bristen på en tydlig jordbrukspolitik i vissa utvecklingsländer ; detta sagt utan att förnärma de skötsamma .
Jag tror att kommissionen kan spela en viktig roll med att hjälpa till att utveckla detta .
Ingen jordbrukare , oavsett var han finns i världen , kommer att producera något om priserna är för låga .
Regeringarna i utvecklingsländerna står alltid inför ett svårt val : vem skall de stödja , jordbrukarna eller människorna i storstäderna som vill ha billiga livsmedel ?
Det gäller att finna denna vanskliga balans tillsammans med kommissionen ; kommissionen skall inte göra det ensam : i de flesta länder där kommissionen är aktiv ger även medlemsstaterna själva utvecklingsbistånd .
Det får inte förekomma att medlemsstaternas politik är raka motsatsen till kommissionens .
Det åvilar kommissionens delegationer att spela en ledande roll vid utvecklingen av den politiska dialogen i utvecklingsländerna och att sörja för att alla länder följer samma linje .
Det krävs också särskild uppmärksamhet för kostnaderna för produktionsmedlen .
Alldeles för ofta delas konstgödsel , djurläkemedel och många andra saker ut gratis till jordbrukarna .
När projektet efter fem år är avslutat är det också slut med den policyn för gratis utdelning .
Jag tror således att kostnadselementet måste utvecklas från början i policyn för alla projekt , och försåvitt jag vet är detta ännu på långa vägar inte alltid fallet .
Slutligen ställer jag mig frågan om inte fonderna skulle kunna utnyttjas litet bättre .
Varje år upptäcker jag i kommissionens och Europeiska utvecklingsfondens budget att de återigen ligger långt efter i fråga om utnyttjandet av fonderna .
Herr talman , herr rådsordförande , herr kommissionär och ärade kolleger !
Egentligen för vi här en debatt bland övertygade , och det är synd .
Vi borde egentligen tala om samstämmighet i utvecklingspolitiken med till exempel Prodi , som redan från början missat en enorm chans .
Han har låtit splittra upp utvecklings- och samarbetspolitiken på tre kommissionärer , vilket i sig är ett framsteg i stället för fyra , det medger jag , men jag vill låta det vara osagt om detta kan garantera en samstämmig politik .
Vi konstaterar också att det fortfarande finns olika generaldirektorat som ibland har att göra med motstridiga förfarande och argument ovanpå denna politik .
Rådsordföranden kom med ett bra förslag , nämligen om att budgetera Europeiska utvecklingsfonden .
Parlamentet skulle naturligtvis verkligen välkomna detta , och om ni skulle kunna genomföra det vore det en stor historisk seger .
Alltsedan Amsterdam står tre begrepp i centrum : integrering , samordning och samstämmighet .
Jag tror inte att det är särskilt mycket som har förverkligats på dessa tre områden ännu .
När man ber om en rapport om framstegen i fråga om samstämmighet kan det inte vara svårt , såvida man inte helt enkelt måste medge att det över huvud taget inte finns något samstämmighet .
Jag skulle hellre se att det kom en rapport om allt det som för närvarande är osammanhängande och att en systematisk strategi utvecklas för att nå fram till en viss samstämmighet , för vi är ännu så länge långt ifrån det .
Det var en sak i rådsordförandens tal som chockerade mig .
Han säger : " Motsättningar i fråga om politik kan leda till balans . "
Det är mycket riktigt så att det som den ena handen ger kan den andra handen ta tillbaka och omvänt .
Detta leder till stagnation och självbedrägeri , och hela globaliseringen har hittills inte lett till något annat än att det visserligen sker förändringar , men att dessa förändringar bara får fattigdomen att öka .
Detta skulle då vara vår prioritet .
Jag vet att vi gör många bra saker , men låt oss börja med det väsentliga .
Herr talman !
Vi har redan konstaterat att det inte föreligger någon rapport från kommissionen , men jag tänker ta upp tre saker i enlighet med de mål som rådet presenterade i sitt yttrande 1997 .
Det första handlar om konfliktlösning .
Jag har under flera år via rådet och kommissionen försökt få reda på varför ingen av institutionerna aktivt deltar och arbetar för konfliktlösning vad gäller det av Marocko ockuperade Västsahara .
FN har en fredsplan .
Vi borde ta detta tillfälle i akt och avsluta den sista koloniala episoden i Afrika .
Jag vill också ta upp migration .
Jag är oroad över de nya bestämmelserna i partnerskapsavtalet med AVS-länderna , som skall kunna göra det lättare att på lösare grunder utvisa invandrare , asylsökande och flyktingar .
Jag vill också verkligen se EU agera som föregångare när det gäller patent på levande organismer .
Vi vet idag att oftare än var fjärde sekund dör någon av hunger .
Tre fjärdedelar av dem är barn under fem år .
Detta beror inte på livsmedelsbrist , utan på det vi har talat mycket om idag , nämligen på den ökande fattigdomen .
Livsmedelsäkerhet och garanti för biologisk mångfald måste gå före kommersiella intressen .
Jag menar att patent på levande organismer enbart syftar till att kontrollera den globala livsmedelsförsörjningen , speciellt i kommersiellt syfte och inte till någonting annat .
Jag vill också i den rapport som jag hoppas kommer från kommissionen se något om kvinnor .
Kvinnor verkar i alla sammanhang , och inte minst i utvecklingspolitiken , vara fullständigt frånvarande , vilket vi ju faktiskt egentligen inte är .
Herr talman !
Den debatt som vi för idag understryker starkt behovet att diskutera utvecklingspolitik i långt vidare termer än genom att bara mäta biståndsflödena .
Biståndsnivån är naturligtvis viktig , och den bör höjas för de rika länderna i sin helhet .
Detta bör ske inte minst för att bekämpa fattigdomen och genom att satsa på kapacitetsutveckling .
Biståndsnivån är emellertid bara ett av många instrument som starkt påverkar de fattiga ländernas utveckling .
En rad kollegor har idag pekat på områden som utöver biståndet är viktiga och där kontraster och motsättningar mellan olika politikområden är väldigt allvarliga .
Det gäller bland annat handelspolitik , jordbrukspolitik och fiskepolitik .
Andra viktiga områden är naturligtvis flödet av privata investeringar , samarbetet kring forskning och teknologi samt hur världssamfundet hanterar och finansierar olika globala problem som rör oss alla .
Dessa problem omfattar klimatfrågor , biodiversitet , hälsofrågor osv .
Detta konstaterande accentueras av globaliseringen , det vill säga den nya ekonomi som växer fram .
I denna ekonomi är sambanden mellan olika politikområden allt starkare .
Vad vi diskuterar här idag är enligt min mening delvis EU : s bidrag till debatten om globaliseringens möjligheter och risker samt om de spelregler som måste finnas för att ge de fattiga länderna en bra chans .
Den redovisning , eller kartläggning som Maij-Weggen har krävt av hur de olika politikområdena går in i varandra och hur motsättningarna ser ut är naturligtvis helt central .
Jag måste fråga mig varför inte mer har gjorts från kommissionens sida .
Kommissionen är ny , man måste ge den tid , men frånvaron av en sådan kartläggning tyder på att det finns starka spänningar inom kommissionen .
Jag kan bara hoppas att Nielsen skall bli framgångsrik i de kommande diskussionerna inom kommissionen .
Utöver denna typ av redovisning skulle jag vilja se en mer positiv analys som skulle kunna vara löpande .
I denna analys skulle man inte bara titta på biståndsflödena utan övergripande på alla olika typer av stödformer och transfereringar som påverkar de fattiga länderna .
Det gäller teknik , handelsfrågor , samarbete på forskningens område osv .
Det skulle vara ett väldigt konstruktivt bidrag till den debatt som vi för .
Slutligen , i punkt 6 i resolutionsförslaget , rekommenderar parlamentet att en arbetsgrupp tillsätts , för att åstadkomma sammanhållning .
Jag tror att det bara är en tillfällighet , men i denna grupp skall naturligtvis miljökommissionären ingå .
Låt oss hoppas att den debatt vi nu för kommer att vara en vattendelare .
Politiken hittills har alltför mycket präglats av att ge med ena handen och ta med den andra .
Det är många som kommer att följa den fortsatta utvecklingen med stort intresse .
Herr talman !
Demonstranterna i Seattle hävdade att frihandeln är dålig för de mindre och de minst utvecklade länderna : de sade att det är någonting som enbart ligger i de rika ländernas egoistiska intressen .
Och ändå kan vi betänka takten för ekonomisk utveckling och takten för minskning av fattigdom i länder som Indien och Tanzania under de 40 eller 50 år som har gått sedan de blev självständiga .
Där resonerade man att protektionism och statliga interventioner skulle bevara arbeten och göra det möjligt för industrin att anpassa sig gradvis och smärtfritt .
Det fungerade inte ; fattigdomen blev värre än någonsin .
Medicinen kanske inte smakar så gott på kort sikt , men om man öppnar upp sin ekonomi för konkurrens , såväl inom landet som internationellt , tvingar det fram ett optimalt utnyttjande av resurserna , och det leder till en högre levnadsstandard och livskvalitet på inte alltför lång sikt .
Är inte det den lärdom som man kan dra av Europeiska unionen själv , särskilt av den inre marknaden ?
Som Nielson sade , utgör den ett fint exempel för de länder och regioner som strävar efter ökat välstånd .
Men det räcker inte med att predika om frihandelns fördelar för utvecklingsländerna .
Vi måste också leva som vi lär och öka vår egen tillgänglighet för importen från dessa länder .
I parlamentets resolution om WTO-förhandlingarna förordas en öppen importpolitik från EU : s sida .
Denna importpolitik skall avlägsna alla återstående importhinder , tullhinder och kvoter och , något som är lika viktigt , icke-tariffiära hinder , som de exempel Maij-Weggen nämnde i sitt tal - om vi avlägsnade dessa hinder , skulle det göra mer än någon summa utvecklingsbistånd för att säkra den ekonomiska utveckling för utvecklingsländerna som både de och vi önskar .
Det är ganska uppenbart att en brist på samstämmighet mellan utvecklingspolitiken och handelspolitiken försvagar våra ansträngningar på utvecklingsområdet , och den minskar säkerligen också utvecklingsländernas politiska aktning för Europa och våra vackra ord .
Herr talman !
Under de senaste dagarna har vi hört vackra ord om behovet av större samstämmighet , samordning och effektivitet i gemenskapens och medlemsstaternas externa biståndsprogram .
Det finns ett relativt litet verksamhetsområde som är enormt synligt för allmänheten och som skulle vara ett avgörande prov på unionens förmåga att matcha ord och handling .
Jag syftar på den fortgående tragedin med antipersonella landminor , som utgör ett hinder för så många utvecklingsprogram , för återuppbyggnader efter konflikter och som förstör livet för många av de mest utsatta människorna i några av världens fattigaste delar , särskilt i utvecklingsländer .
Under de senaste åren har gemenskapen lagt ned omkring 200 miljoner euro på minröjning , hjälp till offer och sammanhörande verksamheter .
Medlemsstaterna har lagt ned liknande summor .
Men det finns fortfarande en enorm ineffektivitet och en brist på vilja att genomföra en strategi som har överkommits med andra medlemmar av det internationella samfundet för att överkomma problemet med antipersonella landminor inom en begränsad tidsrymd .
Nielson identifierade problemen med bristen på samordnade åtgärder och behovet av att bättre komplettera medlemsstaterna .
Detta har man talat om i många år .
Kommissionen måste genomföra interna organisatoriska förändringar , stärka samstämmigheten och effektiviteten för sina åtgärder , och det vore önskvärt om så skedde med en på lämpligt sätt finansierad central enhet med ansvar för minpolitiken .
Den skulle även behöva snabbare kontrakts- och tillämpningsförfaranden samt en utökad flerårig budgetpost och en kraftigt förbättrad förvaltning av sina program .
En lämplig mönstring av minåtgärdsprogrammens effektivitet måste genomföras i vart och ett av de länder som är allvarligt drabbade av landminor .
I mina ögon inbegrips i frågan om landminor så många av de svårigheter avseende organisation , förfaranden , ekonomisk förvaltning och funktionsduglighet som har hemsökt kommissionen och unionen .
Hör dessa hemsökelser till det förflutna , eller kommer vi att finna att Europeiska unionen på detta relativt kompakta och begränsade området fortfarande är oförmögen att uppfylla sina ambitioner ?
Herr talman , kära kolleger !
Kommissionär Nielson , EU-AVS-avtalet är ett viktigt steg till ökad samstämmighet .
Och det är bra att kriterier som mänskliga rättigheter , demokrati , rättsstatlighet , good governance är bättre förankrade i det nya fördraget än tidigare , att tidigare koloniala förbindelser inte längre så mycket får forma den större delen av våra förbindelser , utan att dessa politiska kriterier har fått större tyngd här .
Detta är nämligen förutsättningen för alla typer av utveckling .
Om dessa kriterier inte uppfylls har utvecklingen inte en chans .
Detta , herr Modrow , gäller även Kuba .
Det gläder mig att Kuba närmar sig denna process .
Men först måste det till en och annan förändring på Kuba .
Alla känner vi till rapporterna från Amnesty International .
Att ni som en av kommunismens sista makthavare har en något annorlunda syn på detta än vad stora delar av denna kammare har liksom att ni har vissa problem när det gäller good governance är ju mycket möjligt .
Icke desto mindre är detta ett viktigt kriterium för Europeiska unionen .
Jag vill föra ett ämne på tal .
Vi talar här om samstämmighet .
Många kolleger har gett exempel på i vilken utsträckning de olika momenten inom politiken inte är samstämmiga .
Men som jag ser det behövs det mer samstämmighet även i utvecklingspolitiken som sådan .
Det är inte samstämmigt att samordningen med medlemsstaterna fortfarande inte fungerar , att det i utvecklingsländer delvis genomförs mycket motstridiga projekt av medlemsstater och Europeiska unionen .
Inte heller är det samstämmigt gentemot den europeiska skattebetalaren att driva en utvecklingspolitik som har underställts unionens budget medan Europeiska utvecklingsfonden fortfarande står utanför .
Herr rådsordförande , om ni i framtiden lyckas med att få dessa 13,5 miljarder euro kontrollerade av budgetkontrollutskottet , att underkasta dem mekanismer som OLAF , då tror jag att ni höjer acceptansnivån .
Jag anser att detta borde vara ett krav även för regeringskonferensen , nämligen att förankra Europeiska utvecklingsfonden i Europeiska unionens budget .
Herr talman , mina damer och herrar !
På det hela taget verkar det finnas goda avsikter bakom denna text , men vi har ändå inte röstat för den i utskottet och vi kommer inte heller att rösta för den i plenarkammaren .
Det finns två skäl till detta , vilket för övrigt fick oss att lämna in några ändringsförslag som jag skulle vilja utveckla mycket kort .
För det första vill utskottet för utveckling och samarbete att Europeiska utvecklingsfonden ( EUF ) överförs till gemenskapspelaren , vilket uppenbart är fel väg att gå .
I våra ögon är samarbetet en mellanstatlig verksamhet , och bör så förbli .
I samband med att Europa är i färd med att förbereda en utvidgning skulle ett införlivande av EUF tillåta vissa att med lätthet dölja deras brist på engagemang bakom den mur som utgörs av gemenskapens budget .
Men då räknar man inte med att vi på så sätt kullkastar ett fruktbart och löftesrikt sätt att ansluta våra partner i Syd till vår samarbetspolitik .
Slutligen har kommissionen nyligen , Maes erinrade lämpligt nog om detta , visat vilka svårigheter som uppstår när den i öppenhet skall förvalta de medel som anslagits till programmen för utveckling och humanitärt bistånd .
Man kan fråga sig varför man skulle skapa ytterligare svårigheter .
För det andra är det för oss mycket beklagligt att man i betänkandet av Corrie nämner handels- och samarbetsavtalet med Sydafrika .
När allt kommer omkring är detta avtal ett praktexempel på den amatördiplomati som Europeiska kommissionen ägnar sig åt , och det i allt större utsträckning .
Man kan med bestörtning konstatera att unionen har kunnat förhandla fram ett avtal för sina medlemsstater , där man utan omsvep ger kommissionen fria händer i fråga om en central del .
Det är än mer skandalöst att rådet har låtit detta ske , så att säga " i förbigående " .
I dag befinner vi oss alltså i en absurd situation , som innebär att vi har försatt oss i ett underläge när vi skall förhandla om så pass vitala aspekter som jordbruks- och vinproduktionen , inom ramen för ett avtal som vi redan har undertecknat .
Den del av avtalet som blockerar förhandlingarna skulle kunna leda till att unionen tvingas ersätta producenter för att sluta framställa sherry , portvin ; en hel rad produkter som enligt den internationella handelsrätten är rena piratkopior , och man kan bara föreställa sig de eventuella kostnaderna för ett sådant prejudikat .
Detta är ett bevis , om vi nu behövde få se fler , på att denna omogna diplomati - som inte försvarar något intresse , med undantag för de särintressen som sitter inkilade mellan frihandelns teologi och mer eller mindre vänskapligt sinnade påtryckningsgrupper och icke-statliga organisationer - inte bara är effektiv , utan också farlig .
Slutligen ett par ord om Corriebetänkandets allmänna inriktning .
I dag betraktar teologerna i Genève och Washington den gemensamma församlingen - låt oss inte dölja det - som ett hinder mot en internationell frihandel .
Det här betänkandet erbjöd ett tillfälle att erinra om att vi bör utveckla och stärka vårt samarbete med länderna i Syd , ett originellt och exemplariskt system .
Det var ett tillfälle som inte utnyttjades i Corriebetänkandet , och vi måste mot vår vilja utdela vårt straff för det faktum att betänkandet är bortkastat på denna punkt . .
( PT ) Herr talman !
För att sammanfatta det sagda skulle jag vilja tydliggöra tre viktiga aspekter i den här debatten .
För det första så kan man rent allmänt säga att det som tagits upp i anförandena är idén om att globaliseringen accentuerar den regionala obalansen och de sociala orättvisorna samt ökar fattigdomen , vilket innebär att något måste göras , annars kommer spänningarna att öka och konflikter uppstå som riskerar freden och den internationella stabiliteten .
För det andra så vore det viktigt att i ett sådant perspektiv se utvecklingspolitiken i en annan synvinkel .
Rollen som den som skall rätta till obalans eller minska orättvisor kanske måste omvärderas .
Det var viktigt att Europeiska unionens roll i den internationella utvecklingspolitiken av alla ansågs vara betydelsefull .
Alla var överens om att Europeiska unionen skulle spela en mera aktiv och ledande roll i den internationella utvecklingspolitiken , men för att göra detta måste man stärka samstämmigheten mellan de olika politikområden som konkurrerar om utvecklingsmålen .
Jag tycker också att det i några anföranden framkom väldigt klart att ansvaret för samstämmigheten mellan olika politikområden inom Europeiska unionen varken tillkommer rådet , kommissionen eller parlamentet ensamt .
Tvärtom bör det vara ett samordnat arbete där eftertanke och lagstiftande och institutionella förberedelser sker i kommissionen eller i rådet och ibland till och med i Europaparlamentet , där för övrigt en del ledamöter redan har lagt fram förslag , som till exempel inrättandet av en kontrollmyndighet eller en arbetsgrupp som skall följa olika politikområden när det gäller utvecklingspolitiken .
Avslutningsvis vill jag påpeka att det också är viktigt att notera att vi måste omvärdera utvecklingspolitiken inom ramen för Europeiska unionens politikområden , särskilt beträffande utrikespolitiken , vilket är en av de frågor som portugisiska ordförandeskapet har prioriterat i sitt program .
Vi menar att detta är absolut nödvändigt .
Vi kommer inte att kunna vidta några logiska åtgärder för att uppnå samstämmighet mellan olika politikområden , om vi inte kan ge utvecklingspolitiken de instrument som behövs för fastställandet av de principer och värderingar som ger Europa dess form i det internationella systemet .
Därför måste vi kanske , som jag tidigare nämnde , byta världsbild och lämna den postkoloniala bakom oss och anamma ett mera europeisk sätt att se på utvecklingspolitiken .
Jag menar ( och även andra noterade detta i sina anföranden ) att antagandet av en ny konvention som kan ersätta Lomékonventionen är ett viktigt reforminstrument och ger ny dynamik åt samtalen med denna viktiga grupp av länder i söder i ett läge när det är viktigt att registrera instabiliteten i de internationella förhandlingar som ägde rum under första förhandlingsrundan i Seattle . .
( EN ) Jag har märkt en viss frustration i många av bidragen till denna debatt .
Jag har på kommissionens vägnar gjort ett uttalande , som jag tror erbjuder en användbar bakgrund till denna diskussion .
Vi kommer att lämna mer detaljerat material som hör direkt samman med alla frågorna om samstämmighet .
Denna diskussion är inte ny .
Vi arbetar för närvarande med den i kommissionen , och när arbetet är slutfört , kommer jag att rapportera om det , eftersom det finns många som har frågat om det kommer att vara möjligt att ta del av rapporten om samstämmighet .
Jag hyser inga tvivel om att det som ett resultat av den ökande politiska uppmärksamhet som dessa problem ges - något som tydligt har speglats i debatten i dag - kommer att bli lättare för kommissionen och Generaldirektoratet för bistånd lyfta fram frågan om samstämmighet till förgrunden av vårt verksamhetsprogram .
Detta kräver också att ytterligare nya mekanismer införs i kommissionssystemet , bland vilka mycket väl kan inbegripas , i enlighet med vad som har föreslagits av vissa av de politiska grupperna i parlamentet , inrättande av en speciell intern arbetsgrupp och upprättande av ett slags för samstämmighetsövervakning i kommissionen .
Jag har läst - och hört under debatten - att man ser på samstämmigheten som en slags mirakelmedel som löser alla problem .
Jag tror att det är viktigt att behålla den som en relativt tydligt definierad disciplin för att försöka minska inkonsekvenser där de verkligen existerar , och vi har sannerligen sådana .
Mycket av detta hör samman med faktiska motsättningar mellan sektorintressen i varenda medlemsstat , och , som det mycket uppriktigt har sagts här i kammaren : människor identifierar sig mer eller mindre med sina intressesfärer , och allt detta är berättigat .
Jag skulle emellertid vilja varna mot illusionen att bristen på samstämmighet är en produkt av någon slags mekanisk ofullkomlighet i systemet .
Det finns sådana , men de utgör bara en liten del av vad vi diskuterar .
Den största delen har att göra med välkända etablerade intressekonflikter mellan till exempel könen , och det är detta som är problemet .
Mulder sade att ingen jordbrukare kommer att börja odla någonting om priset är för lågt .
Detta är sant i vår del av världen , men våra partner och biståndsmottagare i Afrika har ett något annorlunda perspektiv .
De odlar inte bara för att försörja sig , utan för att leva , och det är stor skillnad .
Jordbrukande för att försörja den egna familjen grundar sig inte på prisberäkningar , utan på hoppet om regn nästa säsong .
Detta gäller inte för allt jordbruk i utvecklingsländerna , men för den fattigdomsfokusering som vi måste leverera bättre än hittills .
Med det perspektivet är det som jag säger här av stor betydelse .
Andra frågor har tagits upp : boskapsskötsel i Namibia , tomater och mjölkpulver i Karibien .
Vi bör inte vara för masochistiska .
Det finns en gräns för hur användbart det är .
Alla dessa fall kännetecknas av det faktum att man har tagit hand om dem .
Interventionspriser har reglerats , och de problem som vi hade med nötkött i Västfrika och i Namibia löstes faktiskt genom att interventionsstödet minskades .
Detta är reella problem , men de har alla tagits itu med .
Vad beträffar frågan om kakao , choklad : Jag upprepar att de fem procenten har att göra med att skapa en försörjningsgrund i grannländerna .
Vad vi talar om här är de lokala nötterna , som är lika viktiga för de människor som samlar in dem och försörjer sig på dem i Burkina Faso som kokosnötterna är för odlarna i Ghana .
Detta är inget tydligt fall av brist på samstämmighet , det är mer ett fall av konkurrens mellan leverantörer .
Det som togs upp beträffande socker i Karibien är mer komplicerat .
I " Ramen för utomeuropeiska länder och territorier " utgör ansamlingen av vissa av dessa handelsaspekter ett komplicerat problem , men det kan vara så att vad vi talar om här mer handlar om att främja vissa europeiska företags intressen än om att generera inkomster i Karibien .
Hur som helst är detta en fråga som vi just nu arbetar med .
Jag är fast besluten att försöka skapa en balans i alla dessa frågor , och jag kan nämna framgången med avtalet om handelsutveckling och samarbete med Sydafrika .
I all blygsamhet skulle jag vilja hävda att detta är en sak som bevisar att kommissionen är beredd att gå eller flyga den extra milen för att säkerställa samstämmigheten mellan utvecklingssamarbetesaspekten och handelsintresseaspekten .
Vi har sannerligen gjort vårt för att lösa det problemet , och jag hoppas uppriktigt att vi nu kommer att få en mjuklandning och ett fridfullt genomförande av detta avtal under de kommande åren .
Avslutningsvis tackar jag er återigen för denna debatt .
Vi kommer att återkomma med material om dessa frågor , för dessa problem är här för att stanna , på ett eller annat sätt , av den enkla anledningen att utvecklingssamarbete i grund och botten innebär att göra någonting i världen som innebär någonting annat än att bevaka traditionellt definierade handelsintressen etc .
Vi måste förena dessa olika synsätt .
Tack så mycket , kommissionär Nielson .
Härmed meddelar jag att åtta resolutionsförslag har mottagits i enlighet med punkt 2 , artikel 37 i arbetsordningen .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum på torsdag kl .
12.00 .
 
FN : s nästa session om mänskliga rättigheter Nästa punkt på föredragningslistan är rådets uttalande om unionens prioriteringar inför FN : s nästa session om mänskliga rättigheter den 20 mars 2000 .
Herr talman , ärade kollegor !
Europeiska unionen spelade som alla vet en aktiv roll vid 55 : e sessionen om mänskliga rättigheter i Genève i mars / april 1999 .
Resolutioner om de mänskliga rättigheterna i Iran , Irak , de israeliska bosättningarna , Burma , Myanmar , Republiken Kongo och Republiken Sudan lades fram .
Man formulerade också uttalanden för ordförandeskapets räkning om Colombia och Östtimor .
Europeiska unionen lade för första gången fram en resolution om dödsstraffet , vilken rönte stor framgång och fick stå som förebild för arbetet med resolutionen om barnens rätt , ett gemensamt initiativ med en grupp latinamerikanska länder .
Unionen tänker fortsätta att spela sin roll vid den 56 : e sessionen om de mänskliga rättigheterna i Genève i mars / april .
Särskilt så som överenskommet i rådsgruppen " Mänskliga rättigheter " , Särskilt den 9 februari 2000 då Europeiska unionen , enligt överenskommelse i rådet för de mänskliga rättigheterna , ämnar lägga fram resolutionsförslag om de israeliska bosättningarna , om Iran , Irak och Sudan , om Republiken Kongo och Burma Myanmar samt ordförandeskapets förslag till uttalande om Colombia och möjligtvis om Östtimor , eventuellt som ett förslag till uttalande om situationen i ett flertal länder .
Europeiska unionen fortsätter med sina förberedelser inför den 56 : e sessionen om de mänskliga rättigheterna nästa gång gruppen för de mänskliga rättigheterna sammanträder i mars .
I första hand kommer frågan om ett eventuellt resolutionsförslag om dödsstraff att debatteras .
Hittills har gruppen inte kommit överens om vilken strategi man skall använda för detta , i synnerhet när det gäller utformningen av en kompromiss i sista instans som svar på eventuella ändringsförslag i motsatt riktning , inklusive punkt 7 , artikel 2 i FN-stadgan , som tar upp frågan om suveränitet .
Man försökte enas om ett kompromissförslag efter de svårigheter som uppstod under sammanträdessessionen 1999 i tredje kommittén i FN : s generalförsamling när medlemsstaterna inte kunde komma överens om en ändring i Europeiska unionens resolutionsförslag om dödsstraff eftersom man ville införa en hänvisning till artikel 2.7 .
Förra året , under den 55 : e sessionen för de mänskliga rättigheterna , beslutade Förenta staterna som alla vet att lägga fram ett resolutionsförslag om Kina .
Nämnda resolutionsförslag avslogs efter en kinesisk motion om icke intervention .
Europeiska unionens beslut om vilken attityd man skulle inta gentemot Kina i utskottet för mänskliga rättigheter bekräftades av rådet ( allmänna frågor ) den 21 mars 1999 : inga initiativ från Europeiska unionen om Kina , eller resolutionsförslag om Kina skall stödjas , Europeiska unionen skall rösta mot motionen om icke-intervention .
Det stämmer inte att sammanhållningen inom Europeiska unionen hade bevarats om resolutionen hade gått till omröstning .
Amerikas förenta stater lade fram ett resolutionsförslag om Kina under utskottets 56 : e session om de mänskliga rättigheterna och nu försöker man få Europeiska unionen att skriva under .
Kina har reagerat mycket kraftigt på detta .
De kinesiska myndigheterna står nu i begrepp att vidta rättsliga åtgärder i Europeiska unionens länder och institutioner för att få dem att inte stödja det initiativ som Amerikas förenta stater tagit .
Initiativet debatteras i unionen , inget beslut väntas dock inom kort .
Det ligger i Europeiska unionens intresse att hålla alla vägar öppna så länge som möjligt , åtminstone till efter sammanträdet den 25 februari 2000 där dialogen Europeiska unionen-Kina om de mänskliga rättigheterna skall tas upp .
Med tanke på de ändringar som gjorts av utskottet för mänskliga rättigheter så kan man räkna med att omröstningen om icke-interventionsmotionen kommer att avslås .
Därför är det viktigt att länderna inom Europeiska unionen även i år kommer överens om vilken ståndpunkt som skall intas beträffande en eventuell omröstning av resolutionen .
I det här sammanhanget är det viktigt att notera att Europeiska unionen regelbundet motsätter sig Kinas begäran att dialogen om de mänskliga rättigheterna automatiskt utesluter en resolution i utskottet för de mänskliga rättigheterna i Genève .
Det är uppenbart att Europeiska unionen menar att dialogen samtidigt måste ge konkreta resultat inom området , trots att instrumentet i sig är mycket viktigt för att utbyta synpunkter och för att få reda på vad motparten har för åsikter .
När detta inte sker kan en resolution från utskottet för de mänskliga rättigheterna behövas , eventuellt under dialogens fortskridande .
Europeiska unionen påpekar regelbundet för Kina att utskottet för de mänskliga rättigheterna är rätt instans för att ta upp frågor om de mänskliga rättigheterna och att det , oberoende av om initiativet antas eller inte , i alla fall är berättigat ur den synvinkeln .
Nästa dialog om de mänskliga rättigheterna äger rum i Lissabon den 25 februari .
Seminarier om rättsliga frågor och kvinnans rättigheter kommer att inkluderas och företrädare från den akademiska och civila världen kommer att delta .
Nästa seminarium om de mänskliga rättigheterna som anordnas av det portugisiska ordförandeskapet äger rum i maj 2000 .
Kina godkände vid den senaste rundan av dialogen i oktober 1999 Europeiska unionens förslag om tekniskt bistånd för att stödja ratificeringsförfarandet av det internationella avtalet om ekonomiska , sociala och kulturella rättigheter samt det internationella avtalet om Förenta nationernas civila och politiska rättigheter och som den kinesiska regeringen undertecknat .
Just nu debatteras inom Europeiska unionen de frågor som man gärna ser att Kina åtgärdar .
Som grund för den debatten kommer ordförandeskapet att vidarebefordra ett meddelande till de kinesiska myndigheterna om att Europeiska unionen förväntar sig att Kina vidtar åtgärder vid sessionen den 25 februari .
Ordförandeskapet kommer tillika att överlämna en lista till de kinesiska myndigheterna om individuella fall som vi är särskilt oroade över .
Av sammanträdet som ägde rum i Peking i oktober 1999 framgick att Kina är beredd att göra eftergifter i frågor som har att göra med själva dialogen , med dialogens omstrukturering och med debatten om strafflagstiftning ( dödsstraff , utredningshäktning ) .
Däremot viker de sig inte för de frågor som har att göra med enpartisystemet och territoriell integritet .
Europeiska unionens debatter om situationen i Kina , som ett resultat av dialogerna 1999 , fick Europeiska unionen att bestämma sig för att klargöra sin oro över det som sägs om kränkningar av de mänskliga rättigheterna i Kina och de få konkreta mål som uppnåtts med dialogen , låt vara att man erkänner de steg som i rätt riktning på en internationell plan har tagits av Kina .
Vid ett flertal tillfällen påpekade Europeiska unionen för Kina sitt missnöje med resultatet av dialogen , man hoppades på ett bättre resultat även inom känsliga områden .
Man bestämde sig för att fortsätta med dialogen , men på ett effektivare och mera koncentrerat sätt .
Kina gick med på Europeiska unionens förslag om att omstrukturera dialogen , sakkunniga skall oftare användas och banden mellan seminarierna skall bli starkare .
Vid nästa session för de mänskliga rättigheterna kommer man också att debattera rationaliseringen av det egna arbetet .
Den arbetsgrupp som har till uppgift att granska utskottets rutiner har gjort ett gediget arbete .
Man menar att det är absolut nödvändigt att effektivisera de nuvarande rutinerna och göra dem mera precisa , särskilt inom det finansiella området .
Europeiska unionen kommer att motsätta sig alla falska försök att genom omstrukturering av aktiviteterna i utskottet för mänskliga rättigheter försöka ta bort interventionskapaciteten och minimera handlingsramen och den ständiga uppmärksamheten vad gäller respekten för de mänskliga rättigheterna i världen . .
( EN ) Herr talman !
Jag skulle vilja tacka ordförandeskapet för det förberedelsearbete som det har gjort inför Genèvesammanträdet i frågor som rasism , medborgerliga och politiska rättigheter samt rätten till utveckling .
Som ordförandeskapet sade , återstår mycket att göra , trots den förståeliga begäran från parlamentet och många icke-statliga organisationer om att Europeiska unionen borde offentliggöra sin ståndpunkt i god tid före Genèvesammanträdet .
Det är lättare sagt än gjort - vi diskuterar fortfarande några av de svåraste frågorna .
Till exempel diskuteras många av de saker som togs upp i parlamentets resolution , och det är ännu för tidigt att förutsäga utgången i alla fall .
Det är inte överraskande att debatten är utdragen och svår .
Det är inte ett tecken på någon bristande vilja att förbättra de mänskliga rättigheterna , utan vad det antyder är det vanliga intresset för att få vår strategi rätt , så att vi verkligen får fram vad vill säga .
Låt mig spegla detta intresse genom att ta upp tre kontroversiella frågor : dödsstraffet , Kuba och Kina .
Jag skall vara så oförståndig att jag låter en eller två personliga reflektioner smyga sig in i mina anmärkningar .
Vi undersöker för närvarande alternativen och möjligheterna till att lägga fram en resolution om dödsstraffet i FN : s kommission för mänskliga rättigheter .
Detta har alltid varit en fråga som jag personligen har känt oerhört starkt för ; jag har alltid röstat mot dödsstraffet .
Pådriven av Amnesty International med flera , var ett av de första beslut som jag fattade som guvernör i Hong Kong att avskaffa dödsstraffet .
Vi känner till vad som nyligen hände i FN : s generalförsamling .
Vi var tvungna att frysa vår resolution om dödsstraffet eller riskera att en resolution som skulle ha inbegripet helt oacceptabla argument som hävdade att de mänskliga rättigheterna inte är allmänt tillämpliga och giltiga antogs .
New York-scenen skiljer sig från Genève .
Förra årets debatt i New York om suveränitet och humanitär intervention var ett så känsligt ämne att det påverkade alla andra frågor .
Det påverkade utan tvekan debatten om ett moratorium för dödsstraffet .
Debatten i Genève är emellertid mer inriktad på frågor om de mänskliga rättigheterna .
Vi kan därför ha en bättre chans att göra framsteg där .
För det andra , Kuba .
Jag vill ta upp denna fråga rakt på sak , eftersom vi i Europa med orätt kritiseras för att inte ta de mänskliga rättigheterna där på tillräckligt stort allvar .
Vi är utomordentligt bekymrade över åtgärder från den kubanska regeringens sida under det senaste året som ytterligare har inskränkt den personliga friheten , åtgärder som ändringar av strafflagen och av dödsstraffets omfattning .
Vi oroas också av den senaste tidens ökning av antalet politiska arresteringar .
Vi övervakar situationen för de mänskliga rättigheterna med hjälp av rapporter från icke-statliga organisationer och med hjälp av det arbete som utförs av den arbetsgrupp för mänskliga rättigheter som är baserad på EU-ambassader i Havanna .
Vi har regelbundet framfört vår kritik till de kubanska myndigheterna , och detta parlament har gjort detsamma .
Men jag tror inte att det är rätt strategi att isolera Kuba .
Vi vill se ett Kuba med ett rättvist och öppet samhälle , ett Kuba som respekterar marknadens principer , avtalens okränkbarhet och rättsstatsprincipen .
Vi vill uppmuntra en process med en övergång till demokrati och respekt för de mänskliga rättigheterna och de grundläggande friheterna .
Mina åsikter är exakt desamma när det gäller det tredje ämnet som jag vill ta upp , nämligen Kina .
Kort sagt vill jag att vi skall engagera oss i Kinafrågan .
Det skulle vara slappt och kontraproduktivt , liksom förolämpande mot över en femtedel av mänskligheten , att vilja någonting annat .
Jag vill också se ett Kina som genom fridfulla förändringar omvandlas till ett pluralistiskt samhälle i vilket demokratiaktivister och religionsanhängare inte spärras in .
Så , vad bör vi göra ?
Vi bör naturligtvis bedriva en entusiastisk handel med Kina och hoppas att vi kan välkomna Kina in i Världshandelsorganisationen på vettiga villkor .
Det är felaktigt att tala om en Världshandelsorganisation om inte Kina - eller Ryssland , för den delen - ingår .
Men jag anser inte i dag , och jag har heller aldrig ansett , att vår spirande ekonomiska förbindelse med Kina - som Kinas överskott på 25 miljarder euro i handeln med Europeiska unionen till exempel är ett bevis på - bör tysta oss när det gäller Kinas agerande på området för de mänskliga rättigheterna .
I mina ögon är frågan inte huruvida vi bör ta upp frågan om de mänskligheterna i Kina eller inte - vi har skyldighet att göra det och ett berättigat intresse av att göra det - , utan snarare vilket som är det effektivaste sättet att göra det på .
Så , vilken attityd bör vi ha till en Genèveresolution i år ?
Som ordförandeskapet har påpekat , arbetar unionen som helhet med sin ståndpunkt .
Men jag vill verkligen hävda att det finns ett antal faktorer som medlemsstaterna borde ta lämplig hänsyn till .
För det första , samtidigt som det finns personer som ifrågasätter om det gör någon skillnad att lägga fram en Genèveresolution , anser åtskilliga av de mest framstående kinesiska demokratiförespråkarna att det är ett mycket värdefull steg , inte minst med tanke på det budskap som det sänder till folket i Kina .
Det är en punkt som verkligen är värd att beakta .
För det andra måste vi alla ta lämplig hänsyn till vad som faktiskt har ägt rum i Kina under de senaste månaderna , till exempel de hårda domarna mot demokratiförkämpar , arresteringarna av och straffen som nyligen har utmätts för medlemmar av kristna kyrkor samt arresteringarna av och domarna mot Falun Gong-medlemmar .
De kinesiska ledarna känner väl till vår ståndpunkt i alla dessa frågor liksom i frågan om utvecklingen i Tibet .
Vi har gjort våra åsikter mycket tydliga för dem .
På samma gång som vi alla vet att det för många människor i Kina har skett en påtaglig långsiktig förbättring av deras ekonomiska framtidsutsikter och de sociala och ekonomiska friheterna , har bilden också en mörk sida .
Personer som är kritiska till att lägga fram en resolution säger att vi nu åtminstone för en dialog om de mänskliga rättigheterna med Kina .
Det är sant , och det har ett potentiellt värde , fastän jag måste säga - och jag , liksom ordförandeskapet , har sagt det till kinesiska tjänstemän - att vår dialog inte har haft i närheten så mycket innehåll som vi skulle ha velat .
Naturligtvis har dialogen gjort det möjligt för oss att fastställa och genomföra samarbetsprogram i EU : s regi på det människorättsliga och det rättsliga området .
Det är mycket välkommet , och jag tror också att vårt program för offentlig förvaltning i byar bör hjälpa till att främja demokratin på gräsrotsnivå .
Naturligtvis måste varje dialog som är så komplex som dialogen om mänskliga rättigheter vara en långsiktig process , men jag önskar att jag kunde peka på mer påtagliga framsteg .
Nästa dialog , i Lissabon den 25 februari , kommer att bli ett viktigt prov .
Då kommer vi att se huruvida dialogen leder till resultat eller inte .
Avslutningsvis , vilka är de första steg som vi vill se ?
Ja , till exempel skulle vi vilja se Kina gå från att underteckna FN-konventionerna om medborgerliga och politiska rättigheter samt om sociala och kulturella rättigheter till att verkligen ratificera dem .
Jag önskar att vi var närmare det .
Var står vi då i år ?
Jag upprepar att medlemsstaterna måste bestämma sig .
Vad jag hoppas är , för det första , att vi i Europa kommer att anta en gemensam ståndpunkt och hålla fast vi den , att vi inte kommer att tillåta att någonting tas bort , att vår ståndpunkt inte kommer att grundas på självbedrägeri eller svepskäl , att det kommer att vara en gemensam ståndpunkt och en förnuftig ståndpunkt .
Jag vet att det finns människor som säger att vi måste ha ett bättre sätt för att utöva påtryckningar då det gäller de mänskliga rättigheterna än genom att lägga fram resolutioner .
Men om det är sant , måste vi åtminstone vara mer fantasirika och ärliga mot oss själva i vårt sökande efter denna väg framåt .
Om vi skall vila vår ståndpunkt på dialogen om mänskliga rättigheter , måste vi kunna övertala er , de icke-statliga organisationerna och allmänheten i stort att det verkligen leder någonvart .
Det är , enligt min uppfattning , de närmaste veckornas utmaning .
Jag är tacksam mot kammaren för dess engagemang för de mänskliga rättigheterna runt om i världen , särskilt i Kina .
( Applåder ) Tack så mycket , kommissionär Patten .
Jag förklarar debatten om det gemensamma uttalandet om FN : s nästa session om de mänskliga rättigheterna avslutad .
Vi går vidare med omröstningen .
 
Välkomsthälsning Det är med stor glädje jag välkomnar en delegation från Hong Kongs lagstiftande råd till parlamentet .
( Livliga applåder )
 
OMRÖSTNING .
( EN ) Som Wallström förklarade under gårdagens debatt , kan kommissionen godta följande ändringsförslag : ändringsförslagen 1 , 2 , 7 , 8 , 9 , 10 , 11 och 13 .
Kommissionen kan också godta ändringsförslag 4 i princip .
Kommissionen kan inte godta ändringsförslagen 3 , 5 , 6 , 12 , 14 , 18 och 16 .
( Talmannen förklarade den gemensamma ståndpunkten godkänd ( efter dessa ändringar ) . )
Betänkande ( A5-0023 / 2000 ) av Böge för utskottet för jordbruk och landsbygdens utveckling om förslaget till Europaparlamentets och rådets direktiv om ändring av rådets direktiv 91 / 68 / EEG i fråga om skrapie ( KOM ( 1998 ) 623 - C4-0026 / 1999 - 1998 / 0324 ( COD ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Rekommendation ( A5-0008 / 2000 ) av Cederschiöld för utskottet för rättsliga frågor och den inre marknaden om förslaget till rådets beslut om bemyndigande att på Europeiska gemenskapernas vägnar underteckna WIPO-avtalet om upphovsrätt och WIPO-avtalet om utövande konstnärer och ljudupptagningar ( 11221 / 1999 - KOM ( 1998 ) 249 - C5-0222 / 1999 - 1998 / 0141 ( AVC ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Betänkande ( A5-0015 / 2000 ) av Graefe zu Baringdorf för utskottet för jordbruk och landsbygdens utveckling om förslaget till rådets direktiv om ändring av direktiv 70 / 524 / EEG om fodertillsatser ( KOM ( 1999 ) 388 - C5-0134 / 1999 - 1999 / 0168 ( CNS ) ) Före den slutliga omröstningen : .
( DE ) Herr talman , kära kolleger !
Efter denna omröstning vill jag fråga den ansvarige kommissionär Byrne om han nu , efter att ha sett hur brett stödet är här i parlamentet , är beredd att godkänna ändringsförslagen ? .
( EN ) Jag får tyvärr säga att jag tror att den uttänkta ståndpunkt som jag lade fram i går är den korrekta ståndpunkten .
Den heltäckande strategi som kommissionen har för avsikt att anta för denna fråga kommer att föras fram så snart som möjligt enligt artikel 152 , och parlamentet kommer att ha en medbeslutande funktion .
Det är det bästa sättet att ta itu med detta .
Herr talman !
I enlighet med artikel 69.2 yrkar jag på återförvisning till utskottet .
Motiveringen är att detta handlar om tillnärmning av en lagstiftning som har föreslagits av kommissionen .
Vi har accepterat detta men föreslagit ytterligare tillnärmning av lagstiftning som rör detta direktiv , framför allt när det gäller godkännandet av en text - som i sin helhet har godtagits av kommissionen - om användning och märkning av genetiskt modifierade organismer .
Vi anser att detta hör hemma i tillnärmningen vid detta tillfälle , men kommissionen godtar inte detta .
Jag tycker att vi då i enlighet med artikel 69.2 måste försöka få till stånd ett samtal med kommissionen , och därför ber jag kollegerna godkänna återförvisningen .
( Parlamentet beslutade att återförvisa ärendet till det ansvariga utskottet . )
Betänkande ( A5-0034 / 2000 ) av Stenzel för utskottet för sysselsättning och socialfrågor om utkastet till meddelande till medlemsstaterna om fastställande av riktlinjer för program inom gemenskapsinitiativet Equal för vilka medlemsstaterna uppmanas lämna in förslag till stöd ( KOM ( 1999 ) 476 - C5-0260 / 1999 - 1999 / 2186 ( COS ) ) Före omröstningen : Herr talman !
Låt mig offentligen säga fru Stenzel som medlem av ledningen för ÖVP ( Österrikiska folkpartiet ) att många av ledamöterna här är förskräckta över att ni har ingått en koalition med Haider och att vi fördömer detta !
( Applåder från vänster , kommentarer från höger ) föredragande .
( DE ) Bäste herr Cohn-Bendit , ärade parlament !
Jag anser inte att Europaparlamentet är rätta platsen för att göra så massivt intrång i ett lands inrikespolitik , som ni gör !
Jag kan tala för mitt parti , som var en förkämpe för att Österrike blev medlem och anslöt sig till Europeiska unionen .
Som politisk kraft är vi garantin för att Österrike fortsätter att vara förbundet med de europeiska värderingarna .
Jag vägrar låta mig placeras på högerkanten här av inrikes- och partipolitiska skäl !
Detta har ingenting med sanningen att göra , utan det handlar om ren polemik !
Jag tillbakavisar detta med bestämdhet !
( Livliga , ihållande applåder från mitten och höger , protester från vänster )
 
Välkomsthälsning Detta är kanske ett lämpligt tillfälle att välkomna en delegation bestående av fyra ledamöter från det marockanska parlamentet , ledd av Brahim Rachidi , vice talman i representanthuset , vilken har tagit plats på åhörarläktaren .
Vi är hedrade av denna delegations besök , som äger rum kort före ikraftträdandet den 1 mars 2000 av associeringsavtalet mellan Marocko och Europeiska unionen .
I detta historiska ögonblick välkomnar vi denna utveckling för våra förbindelser och utsikterna till närmare band mellan våra två parlament .
Det är i denna anda som delegationen för förbindelserna med Maghrebländerna kommer att besöka Marocko den 20 till 22 mars .
Jag hoppas att delegationen kommer att ha ett utmärkt besök i Strasbourg .
( Livliga applåder ) Herr talman !
Jag vill bara dra nytta av det faktum att ni välkomnar en delegation , för att meddela att även vi i dag önskar välkomna de ansvariga i de österrikiska antirasistiska organisationer som hedrar oss med att besöka parlamentet .
( Applåder ) ( Sammanträdet avbröts kl .
11.50 för ett högtidligt möte med anledning av ett tal av Vaclav Havel , president i Tjeckiska republiken , och återupptogs kl .
12.50 . )
 
OMRÖSTNING ( fortsättning ) Vi skall nu fortsätta med omröstningen av betänkande ( A5-0034 / 2000 ) av Stenzel om Equal-initiativet .
( Parlamentet antog resolutionen . )
Andrabehandlingsrekommendation : ( A5-0027 / 2000 ) av Lienemann för utskottet för miljö , folkhälsa och konsumentfrågor om rådets gemensamma ståndpunkt ( 9085 / 3 / 1999 - C5-0209 / 1999 - 1997 / 0067 ( COD ) ) inför antagandet av Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapsåtgärder på vattenpolitikens område Före omröstningen : .
( EN ) Vad beträffar kommissionens ståndpunkt i fråga om de ändringsförslag som har lagts fram av parlamentet , vill jag bekräfta vad min kollega sade under debatten här i kammaren tisdagen den 15 februari .
Mer bestämt kan kommissionen godta ändringsförslagen 6 , 16 , 21 , 28 , 31 , 33 , 34 , 44 , 45 , 46 , 48 , 52 , 53 , 65 , 67 , 68 , 75 , 76 , 78 , 80 , 84 , 85 , 88 och 102 i sin helhet .
Kommissionen kan delvis godta ändringsförslagen 8 , 18 , 27 , 29 , 42 , 43 , 47 , 54 , 60 , 62 , 93 , 94 , 104 och 105 .
Kommissionen kan i princip godta ändringsförslagen 2 , 3 , 5 , 7 , 10 , 12 , 14 , 17 , 20 , 22 , 24 , 25 , 26 , 30 , 32 , 35 , 36 , 37 , 38 , 50 , 55 , 56 , 57 , 58 , 63 , 69 , 73 , 79 , 86 , 89 , 96 , 99 , 106 och 108 .
Men kommissionen kan inte godta ändringsförslagen 1 , 4 , 9 , 11 , 13 , 15 , 19 , 23 , 39 , 40 , 41 , 49 , 51 , 59 , 61 , 64 , 66 , 70 , 71 , 72 , 74 , 77 , 83 , 87 , 90 , 91 , 92 , 95 , 97 , 98 , 81 ( rev. ) , 100 , 101 , 103 och 107 .
Tack för er uppmärksamhet .
( Talmannen förklarade den gemensamma ståndpunkten antagen ( efter dessa ändringar ) . )
Betänkande ( A5-0033 / 2000 ) av Andersson för utskottet för sysselsättning och socialfrågor om meddelandet från kommissionen om en samordnad strategi för att modernisera social trygghet ( KOM ( 1999 ) 347 - C5-0253 / 1999 - 1999 / 2182 ( COS ) ) ( Parlamentet antog resolutionen . ) Talmannen .
Jag förklarar omröstningen avslutad Röstförklaringar- Betänkande ( A5-0014 / 2000 ) av Lienemann Jag välkomnar kvaliteten på och ambitionen i betänkandet om Life .
Jag vill kort påminna om att Life är ett finansiellt instrument i miljöpolitikens tjänst , såväl inom Europeiska unionen som i tredje land , vare sig det handlar om grannländerna i Medelhavsområdet , länderna kring Östersjön eller de länder som kandiderar för ett EU-medlemskap .
Utskottet för miljö , folkhälsa och konsumentpolitik har lagt fram många ändringsförslag , och de flesta av dem har införlivats i rådets gemensamma ståndpunkt .
Under den tredje etappen ( 2000-2004 ) kommer Life att delas in i tre huvudinriktningar : Life-Natur ( 47 procent av medlen ) , Life-Miljö ( 47 procent ) och Life-Tredje land ( 6 procent ) .
De viktigaste förändringarna är enligt min mening : Life : s bidrag till en hållbar utveckling inom gemenskapen såväl som en utveckling av gemenskapens politik på miljöområdet , bland annat när det gäller att integrera miljöaspekten inom andra politikområden , samt instrumentets bidrag till miljölagstiftningens tillämpning och modernisering , en förbättrad effektivitet , öppenhet och metod för att genomföra Life , liksom en bättre upplysning och information till allmänheten och ett större samarbete mellan förmånstagarna , Life : s mål bör framför allt vara en hållbar utveckling i tätortsområden , genom en nära koppling med pilotprojekt som genomförts inom ramen för Urban-initiativet , som jag har uttalat mig om på annat håll , de permanenta projektens bidrag till varaktiga sociala och ekonomiska aktiviteter och därmed fler arbetstillfällen .
Det som för mig framstår som ytterst viktigt , är att Life-instrumentet skall förbli öppet för de central- och östeuropeiska kandidatländernas deltagande .
Övriga kandidatländer ( t.ex.
Cypern , Turkiet och Malta ) kommer också att kunna delta i Life , när man har slutit relevanta avtal med länderna i fråga .
Svårigheten i förhandlingarna med rådet handlar givetvis om hur stort totalanslaget för Life-programmets tredje etapp ( 2000-2004 ) skall vara .
Kommissionens förslag , som rådet har bekräftat , ligger på 613 miljoner euro , samtidigt som miljöutskottet har gjort bedömningen att budgeten borde omfatta 850 miljoner euro .
Jag stöder föredragandens beslutsamhet .
Det finansiella anslaget har i själva verket inte anpassats sedan programmet tillkom , inte ens då antalet medlemsstater utökades till femton efter EG : s utvidgning .
Antas detta betänkande i plenarkammaren kommer en förlikning att inledas , i enlighet med medbeslutandeförfarandet , så att vi skall kunna lösa frågan om storleken på programmets medel .
Den här typen av förfarande är en vanlig metod , eftersom program och lagar alltför ofta förses med en budget som inte motsvarar ambitionerna !
Betänkande ( A5-0023 / 2000 ) av Böge .
( FR ) Som ledamot av Europaparlamentet och framför allt som medborgare och konsument , gläder jag mig åt Europeiska kommissionens förslag , som markerar ytterligare ett steg mot en bättre livsmedelssäkerhet inom Europeiska unionen .
Det är ett dubbelt förslag : det handlar dels om att ändra rådets direktiv från 1991 om djurhälsovillkor genom att stryka de bestämmelser som rör skrapie hos får , och dels att inrätta en ny förordning om fastställande av bestämmelser för förebyggande och kontroll av viss transmissibel spongiform encefalopati ( TSE ) , eller sjukdomar av BSE-typ som påverkar får och andra djurarter .
Intressant med den nya lagstiftningen är det faktum att man inrättar en specifik rättslig grund för bekämpningen av skrapie hos får .
Detta gläder mig särskilt , eftersom det var ett av våra främsta krav i uppföljningsrapporten om galna ko-krisen .
Med hänsyn till strävan efter samstämmighet verkar det för övrigt nödvändigt att harmonisera de befintliga lagarna om skrapie - som är begränsade till handeln med får och getter - till ett komplett enhetligt system som omfattar de nya reglerna om TSE , som påverkar alla djur i hela Europeiska unionen , regler som är avsedda att förekomma konsumtionen av livsmedel eller djurfoder .
Denna förordning är särskilt välkommen med tanke på att det fortfarande råder tvivel om skrapie hos får .
Vissa vetenskapliga hypoteser stöder det faktum att skrapie skulle ha kunnat utvecklats till BSE bland nötkreatur och således vara källan till BSE-epidemin .
Även om Europaparlamentets och rådets förslag till förordning om förebyggande och kontroll av vissa former av TSE måste preciseras och stärkas , bland annat vad gäller att spåra och bekämpa skrapie , utgör det en märkbar förbättring .
Det är en garanti till de europeiska medborgarna , som upprepade gånger har vittnat om sin oro över EU : s politik på livsmedelsområdet .
Medborgarnas farhågor , förmedlade av Europaparlamentet , har hörsammats .
Debatterna om försiktighetsprincipen , spårbarhet , ansvar och öppenhet har förmått Europeiska kommissionen att presentera en vitbok om livsmedelssäkerhet .
Denna vitbok presenterar flera tankespår och här föreslås bland annat att man skall inrätta en oberoende europeisk livsmedelsmyndighet .
Allt detta är en del av en europeisk strategi för att återvinna konsumenternas förtroende .
Det är vår sak , ansvariga européer , att visa att livsmedelssäkerheten är förenlig med den inre marknaden och varors fria rörlighet !
Betänkande ( A5-0008 / 2000 ) av Cederschiöld Herr talman !
Jag röstade för förslaget om att göra om lagstiftningen som gäller upphovsrätt , eftersom jag anser att detta är ett av de viktigaste områdena för Europaparlamentet .
Jag anser att det som produceras med tankens hjälp är betydligt viktigare än konstruktioner , konkreta produkter , sådant som vi kan se och röra , eftersom tankemöda och forskning , sådant som man inte kan ta på med händerna , ger resultat av stor betydelse som vi inom Europeiska gemenskapen måste stödja mycket aktivare , inte bara genom att skydda patenträttigheterna utan också genom att bevilja lättnader och stöd åt forskare , åt dem som - genom att utnyttja den utbildning de fått - anstränger sig för att ge kommande generationer något ännu viktigare än det vi fått från det förflutna . .
( DA ) Vi är i princip motståndare till att Europeiska gemenskapen ingår avtal om upphovsrätt på medlemsstaternas vägnar .
Vi noterar emellertid att det handlar om gemensam behörighet mellan medlemsstaterna och gemenskapen , och samtidigt bedömer vi att WIPO-avtalet är ett viktigt framsteg för säkerställandet av distributörers och utövande konstnärers rättigheter .
Vi röstar därför för rekommendationen . - ( DE ) Gruppen De gröna / Europeiska fria alliansen har avstått från att rösta i denna fråga eftersom kommissionär Bolkestein under plenardebatten dagen innan inte svarade på någon av mina frågor gällande EU : s anslutning till WIPO-avtalen ( World Intellectual Property Organization ) .
Institutionellt sett har man inte klarat ut vilken roll Europaparlamentet kommer att spela i vidareutvecklingen av WIPO-fördragen .
Dessutom kan man urskilja en tendens att vid internationella ansvarsuppgifter allt oftare utverka en ren EU-behörighet .
När det då inte står klart i vilken utsträckning Europaparlamentet kan komma att delta i beslutsprocesserna inställer sig frågan om legitimering .
Dessutom har begreppet upphovsman inte definierats i fördragen .
Inte heller här har kommissionen svarat på enligt vilken definition man tänker agera samt huruvida man tänker lösa synliga konflikter genom att påtvinga andra sin egen rättsdefinition .
En av de känsligaste punkterna är allmänhetens intresse - kommer införlivandet och tillämpningen av WIPO att leda till privatisering av utbildningen ?
Och slutligen måste frågan om förhållandet mellan TRIPS ( Trade-Related Aspects of Intellectual Property Rights ) och WIPO redas ut - även här endast tystnad som " svar " från kommissionen .
Om en på förhand utlyst parlamentsdebatt inte har någonting att bidra med till ett klarläggande och ståndpunktstagande , då är det minsta vi kan göra att avstå från att rösta !
Betänkande ( A5-0015 / 2000 ) av Graefe zu Baringdorf .
( PT ) Livsmedelssäkerhet är fortfarande en central fråga efter skandalerna med BSE och dioxiderna .
Genetiskt modifierade organismer ( GMO ) är fortfarande osäkra kort vad gäller miljöpåverkan och människors och djurs hälsa .
Försiktighet bör därför råda där vetenskapliga bevis saknas .
Användandet av biotekniken måste studeras mera ingående och inte vara " omslaget " och till salu i några multinationella bolags vinstintresse .
För övrigt har vinstintresset varit drivmotor för de nuvarande livsmedelskriserna .
Det är i den här situationen som föredraganden befinner sig i , det vill säga GMO sätts under samma juridiska tak som djurfoder , men kom ihåg att " dessa bara får godkännas om de är oskadliga för människors hälsa och miljön " .
Beakta dessutom att " genetiskt modifierade tillsatser klart och tydligt skall anges på varje etikett , administrativt dokument eller annan typ av bifogat dokument " .
Detta underlättar en kontroll och spårning av ämnena och garanterar att konsumenten fritt kan välja .
Efter avtalet i Montreal om genetiskt modifierade organismer ( GMO ) är det positivt att föredraganden i sitt betänkande har inkluderat den här problematiken , och det var detta som fick mig att rösta för betänkandet .
Betänkande ( A5-0034 / 2000 ) av Stenzel Herr talman !
Jag skulle mycket kort vilja ge en röstförklaring för PPE-DE-gruppens räkning om Equal-betänkandet .
Vi följde en röstlista som var exakt likadan som den vi hade avtalat med den socialistiska gruppen i förväg .
Den socialistiska gruppen tog tillbaka detta , och därigenom är betänkandet nu inte lika tydligt som det skulle ha varit annars .
Det gav oss anledning att avstå från att rösta .
Vi vill se till att Equal-betänkandet , som är mycket viktigt för såväl flyktingarna som pensionärerna , de handikappade och kvinnorna , helt enkelt går igenom .
Det är beklagligt att förfarandet har lett till att detta får en sådan negativ uppmärksamhet under denna session .
Jag är övertygad om att föredragandens nationalitet har spelat en viss roll , vilket inte borde förekomma i detta parlament .
Det strider egentligen mot de europeiska värdena och helt klart mot de parlamentariska värden som det talas så mycket om i detta parlament .
Detta har varit våra skäl för att avstå från att rösta vid omröstningen om detta betänkande .
Vi vill att Equal går igenom .
Vi är överens om en mycket stor del av det , men vi beklagar förfarandet och framför allt att vissa grupper har missbrukat detta förfarande på ett billigt sätt .
Herr talman !
Det var bland annat i min egenskap av företrädare för Pensionärspartiet i Europaparlamentet som jag avstod från att rösta på Equal-initiativet , för även om det på ett bättre sätt än tidigare inför stödet till projekt som är avsedda att bekämpa diskriminering på grund av ålder , så är det inte tillräckligt skarpt och konkret i det avseendet .
Men jag avstod också av en annan anledning : jag tror stunden är kommen för Europeiska unionens institutioner att sluta experimentera och leta efter bra rutiner för det som vi skall göra och i stället börja ge de europeiska medborgarna konkret information om vad Europa vill att Europa skall vara .
Vi måste vidta konkreta åtgärder och övergå från teori till praktik . .
( DA ) Vi har röstat för betänkandet om meddelandet från kommissionen om riktlinjer för program inom gemenskapsinitiativ ( CIP ) .
I grunden är vi emot denna typ av program och strukturfonder , men eftersom omröstningen endast behandlar hur - och inte om - dessa resurser skall användas , har vi bara tagit ställning till detta .
Vi anser att ett säkerställande av lika möjligheter för de grupper som nämns i betänkandet är viktigt . .
( FR ) Vi har inte röstat emot detta betänkande , med tanke på att den innehåller ett antal rättvisa allmänna principer , till exempel kravet på att bekämpa rasism på arbetsplatsen och att minska bristen på jämställdhet på arbetsmarknaden .
Men vi har inte heller röstat för , eftersom detta stannar vid mycket vaga , för att inte säga fromma önskningar .
I kapitlet om stöd- och utbildningsprojekt för flyktingar , markerar betänkandet dessutom ett steg tillbaka i jämförelse med den ursprungliga texten , eftersom man preciserar att det inte längre är flyktingar som sådana som berörs , utan " flyktingar i enlighet med Genèvekonventionen " .
Denna restriktion är oacceptabel med tanke på att många flyktingar i hela Europa befinner sig i en dramatisk situation : skyddslösa , tvingade att arbeta i hemlighet och att hålla sig gömda , eftersom regeringen och polisen i de stater som påstår sig vara demokratiska förföljer dem .
Den första åtgärden som krävs på det här området är att ge dem som lever under illegala förhållanden lagliga medel att leva ett värdigt liv och att kunna arbeta utan att degraderas till paria och offer för skrupelfria arbetsgivare och en mängd administrativa och polisiära trakasserier , varav den främsta är att ständigt behöva leva i fruktan för utvisning . .
( EN ) Jag röstade för Stenzels betänkande om Equal-initiativet eftersom jag anser att det är viktigt att fortsätta det arbete som påbörjades med de tidigare delarna Now , Horizon , Youthstart och Integra i Adapt- och Employment-initiativen .
De läxor som vi har lärt av dessa verksamheter måste vi bygga vidare på .
Equal står för " jämlikhet " .
Det måste leda till jämlikhet .
Jag välkomnar den föreslagna koncentrationen på att främja nya sätt att bekämpa diskriminering och varje form av ojämlikhet på arbetsmarknaden .
Jag ansluter mig också till önskan om att vi skall avlägsna oss från ett omodernt format och sammanföra partner i sökandet efter nydanande sätt att angripa arbetslösheten .
Flexibilitet är ett nyckelord .
Jag tycker att det är djupt beklagligt att det bara finns begränsade medel tillgängliga för detta initiativ .
Under den senaste programplaneringsperioden fanns 9 procent av strukturfonderna tillgängliga för gemenskapsinitiativ .
Siffran är i dag 5,35 procent .
Detta innebär att medlen måste användas så att de ger maximal effekt , och information om framgångsrika partnerskap måste spridas snabbt och vida omkring .
Utskottet för sysselsättning och socialfrågor antog flera av de ändringsförslag som jag lade fram , i vilka till exempel berördes betoningen på tillgången till startkapital , frågan om hur man skall utnyttja nya företagartillfällen i städer , i samhällen och på landsbygden samt kritiken om att företagen deltog i otillräcklig grad i det tidigare initiativen .
Detta innebar ofta att goda projekt inte ledde till verkliga arbetstillfällen .
De positiva erfarenheterna av små initiativtagares nydanande åtgärder äventyrades av deras avstånd till den politiska processen .
Jag betonade också behovet av förebyggande .
Även arbetsmarknadsparternas inblandning måste belysas .
Det måste finnas flexibilitet , och prioritet måste ges till att minska den administrativa bördan .
Det måste finnas flexibilitet även för länder med små budgetar .
Fastän det finns vissa aspekter i betänkandet som jag tror skulle kunna angripas bättre på ett annat sätt , anser jag på det stora hela att betänkandet erbjuder en flexibel och förnuftig strategi och att det bör stödjas . .
( PT ) Med det gemensamma initiativet Equal vill kommissionen ersätta gemenskapsinitiativen Emprego och Adapt samt andra underprogram inom nämnda område - Now ( nya möjligheter för kvinnorna ) , Horizon ( för handikappade ) , Youthstart ( ungdomar på arbetsmarknaden ) och Integra ( för dem som riskerar utanförskap ) - med den försvårande omständigheten att man kraftig har dragit ned på de planerade anslagen .
Det är alltså med det här initiativet som man ämnar utveckla det som kommissionen menar är de nya metoderna i kampen mot diskriminering och all annan orättvisa på arbetsmarknaden , där grunden är de fyra pelarna i arbetsmarknadspolitiken .
Mycket som skall åstadkommas med så små medel .
För att nå framgång med det nya arbetssättet borde de förslag som kommissionen antog ha varit mindre komplicerade , enklare och mera direkta och icke-statliga organisationer borde ha fått vara med redan från början så att harmoni får råda mellan intresseföreningarna .
Man gjorde inte detta .
Vi hoppas att de åtminstone kommer att gå igenom våra påpekanden på nytt . .
( FR ) Det är lyckosamt att Europaparlamentet fullföljer sina initiativ i fråga om bekämpning av diskriminering och ojämlikhet .
De fyra områden som omfattas av Equal-programmet - anställbarhet , företagaranda , anpassningsförmåga och lika möjligheter för kvinnor och män - tycks vara mycket lämpliga .
Men detta betänkande , som förmodligen motiveras av de allra bästa avsikter , går här och var i en riktning som förefaller ytterst riskfylld , då det tenderar att sudda ut begreppen om medborgarskap och legala förhållanden samt skapa en gemensam rätt utifrån en mängd undantag , som en grundval för gemenskapens reflektionsarbete .
Visserligen kan man inte annat än godkänna beslutet att vidta specifika åtgärder för att utrota alla de former av diskriminering på arbetsmarknaden som kan drabba asylsökande , som definitionsmässigt redan är hårt drabbade av sitt öde , men vi måste ändå hålla oss till en juridisk tolkning av detta begrepp , i klartext : det finns all anledning att hjälpa vederbörligen erkända asylsökande som befinner sig i en legal situation , men det förhåller sig på ett helt annat sätt med de många kategorier som räknas upp i betänkandet - personer vars ärende är under handläggning , flyktingar med tillfälligt skydd eller personer som nekas flyktingstatus och som riskerar att sändas tillbaka - för vilka betänkandet föreskriver ett identiskt stöd .
Men de stödåtgärder som föreskrivs i betänkandet riskerar - eftersom definitionerna är hårfina - olyckligt nog att utsträckas till fler grupper : asylsökande givetvis , men också asylsökande vilkas ärende är under behandling och slutligen asylsökande som nekas flyktingstatus och som hotas av utvisning .
Dessa skall enligt betänkandet kunna dra nytta av detta åtgärdspaket , samtidigt som deras förhållanden borde , åtminstone vad gäller de sistnämnda , undanta dem från en integrationspolitik i en gemenskap som inte betraktar deras närvaro som legitim och regelmässig - för vad är en asylsökande som nekas flyktingstatus och hotas av utvisning , om inte en invandrare som lever under illegala förhållanden ?
En sådan signal skulle , avsiktligt eller ej , starkt uppmuntra invandringen , eftersom en ansökan om asyl , beviljad eller inte , skulle vara tillräckligt för att motivera en hel rad stödåtgärder som syftar till att integrera dem på ett varaktigt sätt i arbetsvärlden , i en allmän miljö präglad av brist och där de som lever under legala förhållanden , den utländska eller den inhemska befolkningen , skoningslöst konfronteras med arbetslöshetsproblemet .
Trots de allmänna riktlinjerna , som man bara kan stämma in i , var det därför inte tänkbart för mig att sluta upp kring ett betänkande som i sig bär på ett frö till ett nytt angrepp på begreppen medborgarskap och republikansk legalitet , begrepp som jag anser vara särskilt viktiga .
Betänkande ( A5-0027 / 2000 ) av Lieneman Herr talman !
Vi minns alla en filmsuccé som hette " Cocoon " , där de gamla , efter att ha druckit en speciell dryck , blev unga igen .
Det är med andra ord av den största betydelse att vi ägnar dricksvattnet den största uppmärksamhet och att vi uppmärksamt studerar och godkänner de förordningar som gäller vattnet .
Därför har jag godkänt det här förslaget , men jag vill också understryka min önskan att man framför allt inriktar sig på att se till att vattnets renhet , i det ögonblick det kommer in i våra hus , är så rent som möjligt .
I det förslag som godkänts kan jag också konstatera att där fattas - men jag litar på ett det rättas till i framtiden - ett stöd till dem som renar vattnet i sitt eget hem , i den egna bostaden . .
( EL ) Trots den relativa förbättring av det ursprungliga förslaget till direktiv om vattenpolitiken som skett i och med införlivandet av vissa av Europaparlamentets ändringsförslag i rådets gemensamma ståndpunkt , förblir direktivet tveksamt .
Frågor av särskild betydelse är följande : De nya vattenindikatorerna måste vara obligatoriska .
Åtgärder måste vidtas för att skydda grundvattnet från föroreningar .
Det måste finnas bestämmelser om rening av förorenat grundvatten .
Utsläppet av de omkring 400 farliga ämnena i vattnet måste förbjudas , för det finns i dag inte någon egentlig kontroll över dessa .
Det är nödvändigt att få fram ett system som gör det möjligt att snabbt fastställa föroreningar i vattnet .
I kostnaderna för vattendistributionen måste även miljökostnaderna för distributionen beaktas .
På samma gång som kostnaden för att leverera vattnet i allmänhet skall speglas i varans pris , måste det finns särskilda undantag för regioner där ihållande och omfattande torka kombineras med en svår socioekonomiska situation ( t.ex. fattiga regioner eller sociala grupper ) .
Direktivet måste genomföras snabbare .
Mina ställningstaganden kan , bortsett från ändringsförslag 76 där jag gjorde fel för min avsikt var att rösta för , illustreras med hjälp av följande berättelse : Presumtivt förslag till miljödirektiv : " Europaparlamentets och rådets direktiv som fastställer medlemsländernas skyldighet att på gator , torg och i trädgårdar i de europeiska städerna vintertid hålla en temperatur som inte understiger arton grader " .
Direktivets huvuddrag : a ) varje stad skall skaffa de energiresurser och tekniska resurser som krävs för att uppfylla detta mål år 2012 ; b ) kostnaderna skall fördelas mellan stadens samtliga invånare och utgöra en del av elkostnaderna .
Åsikt från en ledamot från norra Europa : " Det här direktivet är orättvist , eftersom en invånare i Stockholm exempelvis skulle få betala drygt tvåhundra gånger mer än den som bor i Neapel . "
Åsikt från en ledamot från södra Europa : " Här rör det sig om konkurrenskraft och lika villkor . "
( Slut på berättelsen ) .
Den ledamot som nu motiverar sin röst ser det som positivt att det finns ett gemenskapsdirektiv om vatten , men anser att ett Europa inte kan byggas med hjälp av en miljödogmatism , utan att man gör sig skyldig till en karikatyr av lagen .
Man kan inte behandla länder som drabbas av översvämningar och torka , Medelhavsländerna till exempel , på samma sätt som länderna i norr med riklig nederbörd i form av regn .
Det skulle innebära ett osolidariskt Europa som praktiskt taget omöjliggjorde överledningen av vatten mellan olika magasin i framtiden .
Vi måste än en gång komma ihåg att vi driver ett kontinentalt projekt med en politisk sammanhållning . .
( FR ) Dricka , livnära sig , tvätta sig , odla ... ; vattnet genomströmmar alla våra handlingar i vårt dagliga liv .
Vattnet betraktas med orätt som en oföränderlig och outtömlig resurs , eftersom en så enkel rörelse som att vrida på en kran verkar så självklar .
Men den självklara källan hotar att sina ...
Alla vetenskapliga studier är nu otvetydiga : vattnet kommer att bli den avgörande frågan under de kommande åren , och det redan i morgon .
Men i morgon är det för sent .
Det är i dag dags att klargöra spelreglerna , innan vi alla blir förlorare .
Genom att anta direktivet om vattenpolitiken , onsdagen den 15 februari , bekräftar Europaparlamentet sin ambition att skydda ytvattnet , det marina och territoriella vattnet samt grundvattnet .
Europa förfogar nu över en struktur som gör det möjligt att förhindra en försämrad vattenkvalitet , främja en hållbar vattenanvändning , skydda ekosystemen , bidra till att motverka översvämningar och torka samt eliminera utsläpp av farliga ämnen .
Det är en livboj vi skickar ut - för att rädda vattnet . .
( FR ) Det är med största nöje jag välkomnar detta ambitiösa förslag till ramdirektiv om vatten .
Den miljökatastrof som nu drabbar Donaus flodstränder påminner oss , om det nu skulle behövas , att den mänskliga nonchalansen alltför ofta leder till att naturresurserna äventyras , såsom vattnet .
Syftet med detta förslag till direktiv , som påbörjades 1997 , är att sätta stopp för den hittills fragmenterade lagstiftningen om vatten och att skydda ytvatten , marina och territoriella vatten samt grundvattnet .
Förslaget erbjuder en struktur som gör det möjligt att förhindra ytterligare försämringar , skydda ekosystemen , främja en hållbar vattenanvändning , bidra till att motverka översvämningar och torka samt att gradvis eliminera utsläpp av farliga ämnen .
Mer specifika direktiv kommer så småningom att antas inom ramen för detta förslag till direktiv .
Det har tagit lång tid att utarbeta denna text .
Förslaget till direktiv har ändrats vid två tillfällen , en första gång 1997 och en andra gång 1998 .
I januari 1999 möttes rådets och parlamentets företrädare i en teknisk arbetsgrupp för att söka sammanföra de båda institutionernas ståndpunkter .
Utskottet för miljö , folkhälsa och konsumentfrågor kom trots det att lämna in många ändringsförslag .
Jag stöder flertalet av dem .
När det gäller tidtabell och mål , föreskriver rådet att målet att uppnå en god ytvattenstatus skall förverkligas senast 16 år efter det att direktivet har trätt i kraft - utskottet för miljö , folkhälsa och konsumentfrågor önskar att den tidsfristen kortas ned till 10 år .
Utskottet kräver också att utsläpp och läckage av farliga ämnen skall ha upphört år 2020 .
Det slutliga målet bör vara att år 2020 ha nått värden som gränsar till noll .
Rådet hoppas på att nå en god grundvattenstatus efter en period om 16 år , men kommissionen har för avsikt att stoppa försämringen av den kemiska kvalitativa grundvattenstatusen för att nå en god grundvattenstatus inom tio år .
Alla de normer och mål som avser skyddade områden bör förverkligas inom tio och inte 16 år .
Jag måste säga att jag är positiv till denna snävare tidtabell , eftersom man också har föreskrivit undantag .
När det gäller kostnaderna godtar jag förslaget som innebär att medlemsstaterna senast år 2010 skall se till att prispolitiken för vatten ger tillräckliga incitament för en effektivare användning av vattenresurserna .
På samma sätt förväntar jag mig att Europeiska kommissionen skall göra ett tydligt uttalande och därigenom åta sig att senast år 2012 lägga fram ett förslag i syfte att säkerställa att miljö- och resursförbrukningskostnaderna avspeglas i priset för vattenanvändningen .
Jag skall avsluta genom att citera ett av ändringsförslagen från utskottet för miljö , vilket inte kräver någon kommentar : " Vatten är ingen vara vilken som helst utan ett arv som tillhör Europeiska unionens folk , ett arv som måste skyddas , förvaras och behandlas som ett sådant . " .
( EN ) Jag vill till det officiella protokollet föra mina åsikter om Lienemannsbetänkandet liksom anledningarna till mitt sätt att rösta .
Vi har alla enats om behovet av att få på plats lämpliga kontrollmekanismer för att skydda våra vattentillgångar liksom mekanismer för att kontrollera vattenanvändarna .
Det finns mycket att hylla i det sätt att angripa problemet som föreslås av föredraganden .
Frågan om skatter eller avgifter på vattenanvändning är emellertid en fråga som , enligt subsidaritetsprincipen , bör lämnas till medlemsstaterna att besluta om .
Enligt min åsikt är det felaktigt att använda ett så trubbigt verktyg som en gemensam europeisk avgift i denna fråga .
I Irland betalar redan alla de stora vattenanvändarna - kommersiella , industriella och inom jordbruket - för sin vattenanvändning .
Detta är ett beslut som bör fattas på nationell eller lokal nivå , och det är på den nivån alla framtida beslut bör fattas .
Dessa är de huvudsakliga skälen till mitt sätt att rösta . .
( EN ) Europeiska unionen är för närvarande i färd med att anta en ny vattenlagstiftning för Europeiska unionen för att uppdatera och upprätta en långsiktig strategi som skall säkerställa tillgången på rent dricksvatten och skydda nuvarande vattenresurser , inklusive floder och kustnära vatten .
Jag stöder målen i denna gemenskapsåtgärd på vattenpolitikens område .
Jag stöder emellertid inte förslaget om att de enskilda vattenanvändarna skall påläggas avgifter för det vatten som används .
Vatten , i detta sammanhang , är en kommersiell handelsvara .
Det är en grundförutsättning för livet självt , och människorna måste ha fri tillgång till den mängd vatten som behövs för det dagliga livet . .
( PT ) Det är positivt att man försöker hejda nedsmutsningen av vattendrag , något som är alarmerande och som regeringarna alltför ofta tenderar att försumma .
Alla vet vi att vatten är fundamentalt för mänskligheten och att vi snabbt måste vidta kvalitetsbevarande åtgärder .
Det är dock lika viktigt att ha i åtanke att vattenpolitiken inte går att särskilja och att ett agerande villkorar alla parter .
Nåväl , såväl i debatten som i förslagen prioriterades frågan om " vattnets fysiologiska , kemiska och ekologiska kvalitet " , bara marginellt nämndes andra skadliga effekter .
Därför måste vi beakta medlemsländernas mångfald , klimatologiska olikheter , hydrologiska betingelser och årets förändringar samt de sociala , ekonomiska och ekologiska effekterna av en tillämpning eller icke tillämpning av normerna .
Det var oron över de här frågorna som fick oss att motsätta oss några av de förslag som utskottet för miljö , folkhälsa och konsumentfrågor lade fram , framför allt de som hänvisar till en alltför strikt kalender och där för litet hänsyn tas till de sociala aspekterna och jordbruket , mycket viktiga för ett land som Portugal där vattenbrist är ett faktum och där den socio-ekonomiska utvecklingen fortfarande är otillräcklig .
Vi menar också att kommissionens och rådets förslag många gånger är alltför bakåtverkande , vi försöker därför vara en jämvikt mellan de villkorliga förslag som har lagts fram . .
( FR ) Rådets gemensamma ståndpunkt om detta förslag till ramdirektiv gjorde oss besvikna .
Den innebär ett minimalistiskt förhållningssätt på många punkter , framför allt när det gäller vilken tidpunkt ett stort antal bestämmelser skall träda i kraft samt antalet undantag och villkoren för att tillämpa ett undantag .
Men det största problemet ligger i definitionen av det mål som Europeiska unionen önskar sträva efter med hjälp av denna text .
Målet är givetvis att i första hand skapa en tydlig allmän struktur , som äntligen skall göra det möjligt att förenkla den tillämpliga rätten i frågan .
Men bortsett från detta bör unionen ha ambitionen att förbättra kvaliteten på såväl ytvattnet som grundvattnet .
Det som står på spel är folkhälsan , dricksvattenförsörjningen , den biologiska kvaliteten och mångfalden , bevarandet av landskapen och djur- och växtarter .
Ur den synvinkeln är den gemensamma ståndpunkten svag .
Jag skulle önska att parlamentet försvarade en mer ambitiös ståndpunkt än rådets , men jag skulle också önska att denna ståndpunkt var trovärdig .
Kravet på " noll utsläpp " och " noll föroreningar " , vilket naturligtvis också gäller de ämnen som finns naturligt i vattnet , är inte realistiskt .
Jag tillhör inte de ledamöter som anser det nödvändigt att anta " extremistiska " ändringsförslag vid andra behandlingen , med det enda syftet att skaffa sig ett handlingsutrymme inför utsikten till en förhandling med ministerrådet .
Jag vill tvärtom ifrågasätta denna strategi som nu har blivit systematisk .
Den skadar parlamentet .
Våra budskap till medborgarna och rådet blir diffusa och inte särskilt trovärdiga .
Alltför strikta miljömål som innebär att hänsyn inte tas till verkliga omständigheter kommer inte att tillämpas , eftersom de aldrig kan uppnås .
Är det vårt budskap , som vi vill föra fram ?
I övrigt finns det en punkt som är särskilt viktig för mig : medlemsstaterna bör kunna , när de så önskar , besluta att upprätta transnationella vattennät .
Den typen av projekt uppfyller principen om sammanhållning och regional solidaritet , vilken vi alltid har försvarat .
Ett sådant projekt bör därför kunna få stöd från Europeiska unionen , inom ramen för främjandet av transeuropeiska nät och regionalpolitik ( via strukturfonderna ) .
Jag vill erinra om att kammaren för två år sedan antog ett initiativbetänkande om de hydrauliska transeuropeiska nätens tekniska genomförbarhet , och jag skulle uppskatta om Europeiska kommissionen under den närmaste tiden kunde informera Europaparlamentet om hur den avser att följa upp det betänkandet . .
( ES ) Vi har blivit vittnen till hur ett betänkande som värnar om Europas vattenkvalitet förvandlas till ett instrument i ett handelskrig .
Vi är alla överens om att vattenkvaliteten är att betrakta som ett mycket viktigt mål , särskilt med tanke på de ofördelaktiga konsekvenser som utvecklingen av modellen för en snabb industriell tillväxt har fått för naturen .
Det är uppenbart att resultatet av denna modell i form av privata vinster har varit olycksbringande , och därför är principen om att förorenaren betalar lämplig för att ta itu med de konsekvenserna .
Men bortom dessa principer ligger synen på vattnet som en gemensam resurs som inte kan underkastas marknadens regler .
Något överraskande , och förmodligen med goda intentioner , har det ekologiska målet förvandlats till ett instrument i ett handelskrig genom att konsumenterna , i synnerhet inom jordbrukssektorn , har fått stå för samtliga kostnader i samband med installationerna och standardanpassningen av dessa .
Sanningen är den att vattnet har blivit ytterligare en handelsvara som är underkastad marknadslagarna .
Det innebär en fullbordad tillämpning av den nyliberala modell som härskar på vattenområdet .
När ingen åtskillnad görs mellan länder och regioner där tillgången på vatten är riklig och inte utgör något problem och regioner där torkan och den låga nederbörden förvandlar vattnet till en knapp resurs som omintetgör möjligheterna till minsta ekonomiska och sociala utveckling , då förstörs den ekologiska principen och vattnet förvandlas till ett kastvapen .
På samma sätt är det ganska ironiskt att möjligheterna försvåras att dela denna resurs som det är så ont om i vissa områden , genom att de som bor i regioner med rikligt med vatten råder invånarna i områden med torka att spara på vattnet .
På grund av denna brist på lyhördhet och solidaritet har jag , som ledamot från en av de torra jordbruksområdena vid Medelhavet men med erfarenheter från områden som Murcia , tvingats att rösta i enlighet med denna framställning . .
( EN ) På Europaparlamentets arbetarpartis vägnar vill jag tala om att vi även om vi har stött den största delen av Lienemannbetänkandet har vissa reservationer .
Den tidtabell som föreskrivs i betänkandet , år 2020 , är orealistisk och ogenomförbar , men den tidtabell som rådet ställer upp , år 2034 , är allt för långt fram i tiden .
Vi tror därför att en förlikning kommer att få fram ett mer realistiskt datum .
Vi har röstat mot ändringsförslagen 25 och 72 , som skulle innebära ett krav på att uppnå en minimal antropogenisk förorening i alla grundvatten .
Vi anser att detta krav är orealistiskt med tanke på de mycket höga kostnaderna och den ytterst långa tidsrymd som ett återställande till en standard nära den ursprungliga skulle kräva .
Det ovanstående förklarar vårt sätt att rösta . .
( FR ) Vattnet är en förnybar och begränsad naturresurs .
En god vattenhushållning är avgörande .
Ramdirektivet om vatten kommer att bli en hörnsten för gemenskapens politik på det här området .
Dess mål är tydliga och ambitiösa .
Vi står bakom dem .
Mängden farliga ämnen som tillförs vattenmiljön fastställs till nära noll .
Men vi anser att det vore klokt att inte införa orealistiska tidsfrister , som varken staterna eller industrierna kommer att kunna respektera .
Visst krävs det en tidtabell , men den måste innehålla fler gradvisa steg .
Den legala förpliktelsen att uppnå noll föroreningar och att utsläppen skall upphöra inom 20 år skulle innebära ett förbud mot alla identifierade ämnen .
Sådana bestämmelser riskerar att skapa stora problem för oss när det gäller gränsöverskridande vattenområden , och för kandidatländerna , vilket hotar att försvåra utvidgningen .
Jag skulle - givetvis - vilja tala om en särskild sektor som jag följer på mycket nära håll , nämligen jordbruket , som är en storkonsument av vatten : jordbruket bör , vilket det redan har börjat göra , acceptera att den som förorenar skall betala .
Men vi måste också ta hänsyn till jordbrukets särskilda förhållanden och begränsningar , särskilt i torra regioner .
När det gäller de ändringsförslag som rör radioaktiva ämnen , ställer jag mig självklart positiv till kontroller , men då uppstår frågan om den rättsliga grunden , som lyder under Euratomfördraget .
Betänkande ( A5-0033 / 2000 ) av Andersson EDD-Gruppen har inte kunnat rösta för Anderssonbetänkandet .
Det finns ju vissa vackra formuleringar , bl.a. erkänds på sidan 15 i motiveringen att " medlemsstaternas olika utvecklingsnivåer och traditioner på området social trygghet omöjliggör en enhetlig harmonisering " .
Nu är begreppet " enhetlig harmonisering " ett av dessa tillkrånglade uttryck som fullständigt förvirrar den integrationsprocess det handlar om .
Det är också korrekt , vilket står i motiveringen , att en harmonisering skulle vara skadlig , eftersom " den skulle ställa högre krav på svagare medlemsstater och i likhet med konkurrensen pressa socialt sett mer utvecklade länder till att göra nedskärningar i de sociala trygghetssystemen .
Ingen skulle vinna på en sådan harmonisering " .
Situationen är emellertid den att man upprättar en social modell som i realiteten handlar om en harmonisering , till på köpet en enhetlig harmonisering .
I skäl D betonas att " unionen kan tillföra ett mervärde genom att anta verkliga konvergenskriterier som är bindande och effektiva " , och sedan betonas det i betänkandet att utvecklingen av denna konvergensprocess främjas genom diskussioner mellan Ekofin-rådet och rådet ( arbetsmarknadsfrågor och sociala frågor ) , och slutligen betonar man i punkt 7 att " processen för social konvergens måste åtföljas av en effektiv och ambitiös skattesamordning " .
Här närmar vi oss kärnpunkten i frågan : Detta projekt med den sociala harmoniseringen är inte socialpolitik , det är en uppföljning av EU : s EMU-projekt , som har ett ganska speciellt intresse för de tre länder som står utanför och som kan rädda sig från detta Titanic , dvs .
Storbritannien , Sverige och Danmark , och det är därför viktigt för oss att betona att vi inte kan stödja ett förslag om viktiga underliggande aspekter syftar till att utvidga EMU-projektet .
Herr talman !
Jag röstade för kommissionens meddelande om en modernisering av den sociala tryggheten eftersom förslaget , enligt min mening , har som mål - även om det inte når ända fram - att äntligen kunna erbjuda en europeisk lagstiftning när det gäller sociala frågor och pensioner .
Jag har lyssnat på de tidigare anförandena med en viss bitterhet , även om jag anser att andan i detta betänkande innebär ett försök att ge ett bättre skydd åt de äldre .
Och detta trots att vi vet att regeringarna i de femton medlemsstaterna skulle vilja skära ner pensionerna så mycket det går .
Jag hoppas verkligen att parlamentet snart har en möjlighet att lagstifta när det gäller pensionerna .
De äldre väntar på att Europaparlamentet skall ge dem en möjlighet att leva bra och i värdighet , bättre än de lever för tillfället .
De nationer som är mindre utvecklade måste nå upp till samma nivå som de stater som , inom Europeiska unionen , garanterar ett bättre socialt skydd . .
( DA ) De danska socialdemokraterna i Europaparlamentet har i dag röstat för betänkandet av vår svenske socialdemokratiske kollega Jan Andersson om kommissionens meddelande om en samordnad strategi för att modernisera social trygghet .
Kommissionens meddelande tar sin utgångspunkt i genomförandet av EMU , som med kravet på stabilitet och tillväxt skapar grunden för att medlemsstaterna skall kunna bevara de sociala trygghetssystemen .
Det fastslås i betänkandet att en modernisering inte betyder att det sker en sänkning av nivån i den sociala tryggheten , utan ett bättre utnyttjande av befintliga resurser .
Vi noterar också att det man i motiveringen fastslår att en modernisering inte heller innebär en harmonisering av de sociala trygghetssystemen , och att en harmonisering tydligen skulle vara skadlig , eftersom den skulle ställa större krav på de svagare medlemsstaterna och i likhet med konkurrensen skulle kunna pressa andra till att skära ned .
En situation som ingen skulle vinna på .
Både i meddelandet från kommissionen och i betänkandet från Andersson , betonas att det är medlemsstaterna som har ansvaret och därmed också bestämmer innehållet i de sociala trygghetssystemen .
Samarbete kring dessa frågor i EU-regi skall tillföra ett mervärde som är grundat på utbyte av erfarenheter , ömsesidig bedömning av utvecklingen av politiken i syfte att fastställa bästa metoder . .
Vi anser att betänkandet innehåller många bra praktiska förslag som vi stödjer , men vi är mycket kritiska till det konvergensperspektiv som genomsyrar betänkandet .
Speciellt vänder vi oss emot de avsnitt som handlar om skatteharmonisering och om att kommissionen skall styra medlemsländernas uppförande ( se t.ex. punkt 7 ) .
Vi vill understryka att området social- och trygghetspolitik i huvudsak skall vara medlemsländernas sak , även om utvidgningen av EU kommer att kräva större samordning än tidigare . .
( FR ) De nuvarande problemen i våra sociala trygghetssystem beror framför allt på ett underskott av intäkter , till följd av arbetslöshet , fattigdom och befolkningens åldrande ; det hänger inte samman med alltför stora utgifter .
Europeiska unionen bär för övrigt ett stort ansvar för denna situation , på grund av den politik som har förts .
Visst måste vi anpassa dessa system .
I bland annat Frankrike måste vi sätta stopp för det faktum att det endast är inkomster av arbete som finansierar sjuk- och pensionsförsäkringarna .
Det krävs också en reform av den föråldrade förvaltningsstrukturen , som är en källa till orättvisor , ekonomisk oreda och slöseri .
Man måste framför allt bedriva en familjepolitik för befolkningstillväxt och en ekonomisk , monetär och finansiell politik för att skapa tillväxt och återerövra den inre marknaden , vilket skulle generera arbetstillfällen .
Vad som föreslås av kommissionen och i betänkandet av Andersson är inte en social politik , det är ett medel att ge Bryssel en orimlig beslutsmakt över finansieringen och därmed över organisationen av och ersättningarna inom de sociala trygghetssystemen i Europas nationer .
Därför har vi röstat emot denna text .
Den sociala tryggheten bör i första hand förmedla den nationella solidariteten .
Och denna solidaritet lyder främst och uteslutande under nationalstatens befogenheter .
Det sociala skyddet bör vara grundat på principen om en nationell och gemenskaplig preferens .
I annat fall blir detta skydd endast ett sätt att ekonomiskt hantera de svåra sociala omständigheter som beror på invandringen , på bekostnad av och till nackdel för den europeiska medborgarna . .
Vi har avstått från att rösta om Jan Anderssons betänkande om en samordnad strategi för att modernisera social trygghet .
Vi har en positiv grundinställning till Europeiska unionen .
Som svenska liberaler ser vi den europeiska integrationen som en möjlighet att nå lösningar på gränsöverskridande problem , såsom miljö , handel , rörlighet över gränserna , mänskliga rättigheter och konflikthantering. gäller det har Europas demokratier en chans att visa världen att samarbete leder till fred och ökat välstånd .
Vi tror också på subsidiaritetsprincipen , att beslut skall fattas så nära den det berör som möjligt .
Det är därför vi aktivt driver frågan om en konstitution för Europeiska unionen , där ansvarsfördelningen är tydlig för envar .
Det måste stå fullkomligt klart för alla medborgare att EU enbart skall syssla med de frågor man kan bäst - de gränsöverskridande .
Alla andra frågor bör hanteras på lokal , regional eller nationell nivå .
Socialpolitik är ett exempel på ett område där EU bara bör ha begränsad kompetens , förutom då det berör den fria rörligheten för människor inom unionen .
Varje medlemsstat bör ha det fulla ansvaret och rätten att själv besluta om sina sociala trygghetssystem .
Sjukvård , barnomsorg och äldreomsorg är tydliga exempel på områden som inte är direkt gränsöverskridande .
Detsamma gäller arbetsmarknadspolitiken .
Vi tror inte att en gemensam europeisk lagstiftning på dessa områden är en lösning på trygghetssystemens problem .
För oss är det viktigt att EU i stället koncentrerar sig på ett fåtal områden där man verkligen kan göra nytta .
Det hindrar däremot inte att medlemsländerna samarbetar och utbyter idéer på det sociala området .
Trygghetsfrågor och jämställdhet är frågor som traditionellt står högt upp på vår liberala agenda .
Flera av de idéer som presenteras i Anderssons betänkande sluter vi helhjärtat upp bakom på nationell nivå . - ( IT ) Vi ser med intresse och förhoppningar fram emot en samlad strategi för att modernisera de sociala trygghetssystemen i Europa , något som emellertid inte får genomföras isolerat från sammanhållningsprocessen : en modernisering , men samtidigt en sammanhållning - detta är något som framkommer i föredragandens betänkande och som vi instämmer i .
Många politiska program har redan , även om det skett med viss möda , slagit in på denna väg , men många andra måste fortfarande göra det innan Europa , även om det bara gäller subsidiariteten , verkligen är ett gemensamt hus , inte bara för medborgarna i medlemsstaterna , utan också för medborgarna i kandidatländerna .
De sociala trygghetssystemen i Europa har för övrigt dessutom alltid spelat en positiv roll när det gäller den civila och demokratiska utvecklingen för Europas folk .
Och om de systemen i dag , med den utveckling som sker inom ekonomi , arbetsmarknad och samhällets behov skall kunna fortsätta vara ett stöd för utvecklingen , så krävs det utan tvekan en modernisering .
De aspekter som vi emellertid måste understryka , är tre : den första gäller det nära inbördes beroende som måste finnas mellan ekonomisk politik , arbete och social trygghet i strikt proportionella termer .
Den andra gäller administrationen av de sociala trygghetssystemen och de organ som ombesörjer detta .
Allt oftare och allt effektivare arbetar man i själva verket i dag med kompletterande och integrerade stödsystem .
Men det som , enligt vår mening , inte kan skäras ner är de offentliga institutionernas roll , såväl vad gäller universaliteten som - hoppas vi - kvaliteten när det gäller att tillhandahålla den sociala grundtryggheten .
Detta är , i allt väsentligt , en fråga om rättvisa och gäller sjukvården , pensionerna och även de fall där det krävs en strategisk samordning , och förnyelse , av den offentliga myndigheten .
Den tredje aspekten gäller subsidiaritetsprincipen , som Europa vilar på .
Det saknas fortfarande en gemensam strategi för det sociala skyddet och den sociala tryggheten , och de system som finns baseras i huvudsak på de åtgärder och den solidaritet som visas inom varje medlemsstat .
En moderniseringsprocess när det gäller de systemen kan inte ignorera skillnaderna vad gäller ekonomi , sysselsättning eller social trygghet mellan de enskilda staterna , oavsett om de är medlemmar eller kandidatländer .
Det krävs med andra ord att moderniseringen , som är nära knuten till en samordningsprocess även om den har olika utgångspunkter , vill och kan inleda en positiv utveckling och inte tvärtom .
Det handlar dessutom om kultur , om framsteg och värdighet i den nuvarande Europeiska unionen och i en framtida utvidgad union . .
Den värdegrund som är gemensam för medlemsländerna i Europeiska unionen bygger på demokrati , mänskliga fri- och rättigheter samt en social marknadsekonomi .
Dessa värderingar måste ges uttryck i solidariteten med de svagare grupperna i vårt samhälle och i omvärlden .
I enlighet med subsidiaritetsprincipen är det medlemsländerna som själva utformar sina sociala trygghetssystem .
Dock bör invånarna i Europeiska unionens länder kunna åtnjuta ett minsta sociala skyddsnät oavsett i vilket land de bor .
I betänkandet efterlyses en " effektiv och ambitiös skattesamordning " utan att närmare definiera innebörden .
Ett sådant ställningstagande är enligt vårt synsätt ett alltför stort ingrepp i den nationella skattepolitiken och kan därför inte stödjas .
Därmed röstar vi emot punkt 7 i betänkandet .
I betänkandet betonas den sociala dimensionen i det europeiska samarbetet , vilket välkomnas .
Det är dock viktigt att klargöra vilken roll EU skall spela , och inte spela , beträffande social trygghet .
Ett sådant klargörande saknas i betänkandet , vilket är beklagligt . .
( EL ) När man läser det av si och så många goda föresatser genomsyrade meddelandet från kommissionen om social trygghet , frågar man sig om de personer som sammanställt meddelandet och de europeiska arbetstagarna lever på samma kontinent , i samma sociala verklighet .
Man frågar sig också om denna " samordnade moderniseringsstrategi " inte är en annan falsk benämning på det samordnade frontalangreppet på socialskyddet och den sociala tryggheten och på de rättigheter som arbetstagarna har uppnått .
Vi delar ganska många av föredragandens åsikter , men vi delar inte alls hans optimism om kommissionens och rådets föresatser och planer vad den sociala tryggheten beträffar .
De allmänna riktlinjerna för den gällande ekonomiska politiken - stabilitetspakten - och de hårda konvergensprogrammen , som drabbar sysselsättningen hårt och som främjar anställbarheten och en uppmjukningen av den sociala dialogen och arbetsorganiseringen , kommissionens och Europeiska centralbankens beslut om återhållsamma löneökningar , liksom framhärdandet i en sträng finansiell disciplin och en till varje pris säkerställd penningpolitisk stabilitet , tillåter oss inte att hysa några tvivel om målen och avsikterna med den nya strategin .
Dess enda syfte är att jämna vägen och skapa förutsättningar för minskade offentliga utgifter för de sociala skyddsnäten och att mjuka upp själva den sociala tryggheten .
När den sociala tryggheten gång på gång och av många ledare beskrivs som en " kostnad " och ett " hinder " för ökad konkurrenskraft , och när man söker efter metoder att flytta över denna kostnad från företagen till arbetstagarna - - hela tiden , naturligtvis , under förevändningen att vilja skapa arbetstillfällen - - skulle vi förvånas om den nuvarande modellen med en otyglad marknadsekonomi , med ett strikt ekonomiskt synsätt i alla lägen , den av de monopoliska intressena fullständigt beroende , skulle ta medborgarnas grundläggande rättighet till social trygghet och vård under sitt beskydd .
Det är uppenbart att vad som eftersträvas är en överflyttning från de organiserade sociala trygghetssystemen - , som ligger under statlig kontroll , - till privata aktörers trygghetssystem , något som kommer att ge nya vinster till kapitalet och ytterligare tynga ned arbetstagarna , som förutom den högre kostnaden kommer att " åtnjuta " allt sämre sociala tjänster .
Den nya omoraliska konkurrensen mellan de offentliga och privata sociala trygghetssystemen , liksom mellan medlemsstaternas system , utgör inte bara inte en satsning , utan den uppenbarar tvärtom de politiska avsikterna och det outhärdliga tryck som man utsätter de sociala trygghetssystemen för i syfte att nedmontera eller bryta upp dem , till fördel för den privata sektorn och lagen om maximal vinst .
Det är känt att sysselsättningsnivån och sysselsättningskvaliteten även bestämmer kvaliteten på de sociala trygghetssystemen .
Hur kan vi tala om sunda och ekonomiskt hållbara sociala trygghetssystem , när vi framför våra ögon har de miljontals arbetslösa , de fattiga , de marginaliserade , deltidsarbetandets " fattiga arbetstagare " , de från de gällande arbetstidsreglerna undantagna ?
Den sociala tryggheten och socialskyddet utgör en av de europeiska arbetstagarnas största landvinningar , och den kunde göras efter mångåriga strider mot storkapitalets strävanden och med den ständiga solidaritet som är ett kännetecken för arbetstagarna .
I dag i arbetslöshetens och undersysselsättningens Europa är det av högsta vikt att säkerställa en bredare social trygghet och en utvidgning av arbetstagarnas rättigheter , vilket emellertid kräver ett annat system för den ekonomiska och sociala utvecklingen , något som EU , på grund av sin natur och karaktär , inte kan erbjuda .
På grundval av dessa värderingar , vill vi uttrycka vårt kategoriska motstånd mot den " modernisering " av det sociala trygghetssystemet som kommissionen föreslår med sitt meddelande och påpeka att vi inte kan rösta för detta betänkande från utskottet för sysselsättning och socialfrågor .
Jag förklarar röstförklaringarna avslutade .
( Sammanträdet avbröts kl .
13.55 och återupptogs kl .
15.00 . )
 
FN : s nästa session om mänskliga rättigheter ( fortsättning ) Nästa punkt på föredragningslistan är debatten om rådets uttalande om unionens prioriteringar för nästa sammanträde för mänskliga rättigheter i FN ( 20 mars 2000 ) , inklusive situationen i Kina .
Herr talman !
Det är verkligen beklagansvärt att rådets tjänstgörande ordförandeskap inte är närvarande ; det handlar om rådets uttalande och jag tror att det skulle ha varit värdefullt om rådet hade varit här under debattens gång .
Jag vill , för jag tror inte att det är bortkastat , påminna om att det faktum att frågan finns upptagen på föredragningslistan visar på ett behov som alla politiska grupper har uttalat , nämligen att parlamentet håller en debatt inför nästa sammanträde i Förenta nationernas kommitté för de mänskliga rättigheterna i Genève , för att kunna göra sig hörd i en fråga som är så pass känslig och angelägen för parlamentet .
Efter det tjänstgörande ordförandeskapets uttalande i rådet och i kommissionen tror jag att vi alla kan vara överens om att den nuvarande situationen för de mänskliga rättigheterna är långt ifrån den vi alla skulle önska .
Vi kan på unionsnivå inte nog påpeka att situationen inte är helt tillfredsställande , till exempel för även om konventionen om skydd för mänskliga rättigheter och grundläggande friheter är ett vanligt inslag i medlemsstaterna , har inte samtliga stater ratificerat eller undertecknat de därpå följande protokollen .
Dessutom är det en klar nackdel i den här frågan om inte Europeiska unionen undertecknar den europeiska konventionen om skydd för mänskliga rättigheter och grundläggande friheter , med alla de nackdelar som en sådan situation innebär .
Jag hoppas att dessa problem tas upp och behandlas inom ramen för de diskussioner som för närvarande pågår om Europeiska unionens stadga för de grundläggande rättigheterna .
På utrikesnivå anser jag att de punkter vi har tagit med i resolutionen ger oss en vision som påminner mycket om verkligheten och inte väcker någon optimism , herr talman , med tanke på att aspekter som upphävandet av dödsstraffet , den tortyr som fortfarande utövas i många till synes demokratiska länder eller situationen för minoritetsbefolkningar på många ställen på vår jord kräver ett tydligt , synligt och verkningsfullt besked från Europeiska unionen .
Jag anser att resolutionen innehåller en rad viktiga frågor , men jag kommer att uppehålla mig vid en mycket speciell fråga , nämligen behovet av en bättre samordning mellan Europeiska unionen och Förenta nationerna .
Herr talman , i en värld som denna , som allt mer domineras av fenomenet globalisering , inte bara på det ekonomiska området , måste vi ge enhetliga och samordnade besked för att de skall vara verkningsfulla .
För att uppnå en sådan verkan i vårt agerande är det nödvändigt att i praktiken skapa den samordning som saknas i dag .
Därför försvarar parlamentet den nödvändiga principen om att delta i kommittén för mänskliga rättigheter och i andra internationella forum där dessa frågor tas upp och , herr tjänstgörande rådsordförande , parlamentet skulle så snart som möjligt vilja delta i den typen av sammankomster .
Europeiska kommissionen planerar att inom kort , i maj månad , lägga fram ett meddelande om utvecklingen av de mänskliga rättigheternas och demokratiseringens roll i unionens utrikesförbindelser .
Jag vill passa på att uppmana kommissionen att ta hänsyn till det behov av samordning som jag just har påtalat och att man söker nya metoder som stärker den roll som Europeiska unionen , och då särskilt parlamentet , har på området mänskliga rättigheter , i synnerhet ur en samordningsaspekt , genom att ge sitt erkännande av den goda viljan hos de tredje länder som godkänner klausulen om demokrati .
Jag anser att det bör gälla samtliga effekter - och då syftar jag särskilt på budgeteffekten .
Slutligen vill jag även nämna de viktigaste bidrag som det civila samhället kan göra på området , liksom den så ofta underskattade rollen hos de många icke-statliga organisationer som agerar i frågan .
Unionen bör bemöda sig om att erbjuda dem allt det stöd de behöver för att kunna uträtta sitt viktiga arbete .
Herr talman , herrar kommissionärer !
När denna kammare skall diskutera mänskliga rättigheter så löper vi en allvarlig risk att problemen , om man säger så , ytterligare understryks av det klimat i vilket vi uppmanas att diskutera denna så viktiga fråga .
Frånvaron av rådets medlemmar och praktiskt taget samtliga parlamentsledamöter gör att vi inser hur långt det fortfarande är mellan de ädla förklaringarna , högstämda och formellt användbara , och de konkreta handlingarna i det dagliga politiska livet när det gäller frågan om mänskliga rättigheter .
Jag anser att detta parlament , med början från det bidrag som Europeiska unionen kommer att ge till mötet i Genève , har som uppgift att fylla igen detta tomrum och lämna ett bidrag , inte bara när det gäller att göra principförklaringar , utan också när det gäller verkligheten och kanske också lojaliteten .
De mänskliga rättigheterna måste komma loss från en tolkning som enbart är knuten till det ögonblick när de formuleras eller när bestraffningar utdelas .
Vi , i egenskap av Europaparlament , har framför allt till uppgift att förvalta de mänskliga rättigheterna i preventivt syfte .
I det avseendet måste vi kunna exportera en kultur av legalitet , en rättskultur , en rutin när det gäller rättsuppfattningen .
Jag tror att vi definitivt kan se slutet på en lång säsong under vilken fördrag lagts till fördrag och namnteckning till namnteckning .
I dag finns det många , kanske för många , fördrag inom området mänskliga rättigheter : om de fördragen även i fortsättningen enbart skall vara tomma förklaringar så förblir de bara samlingsplatser för onödiga tankar .
I dag måste vi gå vidare till nästa fas i utvecklingen , och det är att dagligen och konsekvent tillämpa det som står skrivet i våra fördrag , även om vi inte får glömma att vissa grundläggande fördrag fortfarande inte har antagits : jag tänker på Romkonferensen och det faktum att 14 av 15 länder i unionen ännu inte har ratificerat fördraget om en internationell brottmålsdomstol .
Jag anser att vi måste utvärdera och ändra vissa av de politiska instrument vi utgår från när vi mäter kvaliteten på de mänskliga rättigheterna på vår planet .
Vi har ofta utnyttjat instrument som , formellt sätt , kan verka betryggande men som , när det gäller politiska resultat , är fullständigt verkningslösa : jag tänker på bruket och ofta missbruket av att införa embargo under de senaste åren och den alltför försiktiga tillämpningen av klausulen om upphävande av avtalen mellan Europeiska unionen och tredje land om det i ett sådant land skulle förekomma kränkningar av de mänskliga rättigheterna .
Jag tror att vi framför allt måste ändra omfattningen när det gäller vår skyldighet att skydda de mänskliga rättigheterna .
Globaliseringen riskerar att få en rent negativ tolkning .
I detta ögonblick ifrågasätts i många länder principen om de mänskliga rättigheternas universalitet .
Man hävdar att många mänskliga rättigheter och rätten till liv som förnekas genom dödsstraffet skulle vara beroende variabler , medan globaliseringen , som ofta ses som något negativt , snarare kan bli det nät som håller samman rättigheter , åtgärder och politik i samtliga länder .
Vi måste med andra ord uppdatera vår aktionsradie när det gäller ansträngningarna att skydda de mänskliga rättigheterna : jag tänker på de sociala rättigheterna , de anställdas rättigheter , arbetslivets kvalitet , nödvändigheten av att kräva respekt för alla de viktiga kriterier som Internationella arbetsorganisationen ( ILO ) angivit .
Jag tänker på rätten till tolerans , rätten till respekt , något som är en rättighet för alla minoriteter , framför allt inom Europeiska unionen .
Jag tänker också på rätten till utveckling , vilket är en folkens rättighet , de folk som i sin tur är summan av alla enskilda individer och varje enskild individ i det folk i vilket vederbörande ingår har rätt till utveckling , en framtid som framför allt skall vara en plats för framtidshopp och tillväxt .
Jag menar att allt detta ingår i ett resonemang , en debatt , ett bidrag som Europeiska unionen skall ge när det gäller frågan om mänskliga rättigheter .
Jag hoppas att Europaparlamentets deltagande i det möte som äger rum i Genève inte bara blir en formalitet , och att det inte bara blir ett tillfälle att lyssna och att berätta utan att det framför allt blir ett tillfälle att bekräfta att frågan om de mänskliga rättigheterna för oss är en central dimension , något som Europeiska unionens , den europeiska nationens , identitet är beroende av och att vi också hävdar de mänskliga rättigheternas universella karaktär , en karaktär som sträcker sig bortom tid och rum .
Vi hoppas att det blir så , och detta är den uppmaning som vi riktar till våra regeringar , inte bara som en ren formalitet .
Herr talman !
Även om kammaren för tillfället är ganska tom så har parlamentet en mycket hög profil inom området mänskliga rättigheter .
Från denna kammare har vi uttryckt vår oro och fördömt regimer som förtrycker , torterar , avrättar och diskriminerar sina medborgare .
Detta engagemang skapar oro och ger effekt .
Det har vi flera gånger sett bevis på .
För två veckor sedan fick jag ett brev från Kinas ambassad i Bryssel .
De uttryckte sin bestörtning över att vi i parlamentet har fördömt Kina och ägnade tio sidor åt att förklara att vår kritik bygger på missförstånd .
Detta brev är bara ett exempel som visar att det vi gör inte klingar ohört , utan att det följs med stor uppmärksamhet av omvärlden .
Detta är bra och visar på den viktiga opinionsbildande roll som Europaparlamentet har .
EU : s roll är viktig.Därför måste vi ha en konsekvent , tydlig och sammanhållen politik inom mänskliga rättigheter .
Nu finns det , trots brevet från Kinas ambassad , verkligen skäl att oroa sig för utvecklingen i Kina .
Denna fråga kommer tillsammans med många andra att diskuteras på mötet i Genève om ett par veckor .
Från den liberala gruppen är vi oerhört angelägna om att EU håller fanan högt och agerar kraftigt vid detta tillfälle .
Jag blev glad när jag hörde kommissionär Pattens inlägg om Kina , men lite oroad när jag hörde rådsordförandens tvekan .
En stark resolution om Kina skulle vara en viktig markering mot ett land där det förekommer systematiska brott mot mänskliga rättigheter .
Medlemmar från den andliga , helt fredliga , men nu förbjudna rörelsen Falun Gong , har återigen utsatts för massarresteringar .
Uppgifter kommer om tortyr , isolering och till och med avrättning .
Årslånga fängelsedomar utdelas utan rättegång .
Hundratals gruppmedlemmar skickas till läger för omprogrammering .
Detta är helt oacceptabelt .
Trakasserier förekommer också mot andra grupper såsom protestanter och katoliker .
Kina påstår sig respektera religionsfriheten , men alltför många fall av våld och trakasserier mot religiösa ledare tyder på motsatsen .
Inte heller finns det några tecken på att situationen i Tibet förbättras .
Därifrån kommer fortfarande larmrapporter om tortyr , fängslanden och trakasserier .
Grundläggande rättigheter accepteras inte i Kina .
Det gör inte heller yttrandefrihet , mötesfrihet och organisationsfrihet .
Nu är inte heller informationen fri .
Kina har de senaste veckorna gjort allt för att strypa tillgången till Internet och för att hindra medborgarna från att kommunicera och få information från andra länder via Internet och e-mail .
Allt detta visar att situationen är bekymmersam , och det finns förstås flera strategier för att agera .
Bilaterala dialoger är ett sätt , men det räcker inte .
Man får inte låta sig luras av att Kina fem i tolv gör en symbolisk handling för att ge sken av att det sker förbättringar .
Mötet i Genève är ett viktigt tillfälle för omvärlden att tala om för Kina att systematiska kränkningar av mänskliga rättigheter inte är acceptabla .
Herr talman !
Till detta parlaments räddande verksamhet hör att man bedriver en konsekvent och aktiv människorättspolitik , håller fanan högt som Malmström uttryckte det .
Samtidigt blundar vi emellertid för unionens egna problem : våld , ojämlikhet , fjärde världens verklighet som en del av EU : s vardag .
Det är alldeles riktigt att vi fäster seriös uppmärksamhet vid de kränkningar av de mänskliga rättigheterna som kommer att diskuteras i Genève .
Den retorik som vi använder oss av har dock ofta inslag av självbelåtenhet som ligger hisnande nära den nordamerikanska människorättsnarcissismen .
Det är direkt skenheligt att fördöma även de grövsta brotten mot de mänskliga rättigheterna i tredje land om vi inte är beredda att sträcka ut en hjälpande hand till verkliga flyktingar och asylsökande , vilkas situation nu håller på att försvåras i Europeiska unionen .
Jag vill i synnerhet fästa er uppmärksamhet på bestämmelser om återtagande , re-admission clauses , som äventyrar Genèvekonventionen och som man borde avvärja .
Om vi inte kan upprätthålla den här höga människorättsnivån för asylsökande har vi inte gjort oss förtjänta av de europeiska värden som enligt Vaclav Havel , som talade här i dag , bildar den europeiska identiteten och av vilka han särskilt lyfte fram respekten för de mänskliga rättigheterna och solidariteten .
Jag arbetade under flera år i Sydafrikas sannings- och försoningskommission , och det var frapperande att se hur en nation under svåra förhållanden strävade efter ett pluralistiskt demokratiskt samhälle av en mer öppen europeisk typ .
Jag befarar att vi nu är på väg i motsatt riktning , mot europeisk slutenhet och apartheid .
Herr talman , herr kommissionär , herr rådsordförande !
Den fråga som det här året bör ställas i Genève , det är med all säkerhet inte frågan om dödsstraffet .
Vi har redan fått igenom tre resolutioner i Genève som avser dödsstraffet .
Men i generalförsamlingen förra året misslyckades vi på grund av ett vilseledande svepskäl , artikel 2.7 , som vi för övrigt har antagit för alla andra texter utan problem .
Frågan om dödsstraffet skall alltså upp i generalförsamlingen i år , och inte vid sessionen i Genève .
Den absolut avgörande punkten , vilken Patten pekade på - och jag vill tacka honom för de ståndpunkter han försvarade - det är Kina .
Tyvärr är avståndet mellan rådets och kommissionens ståndpunkter längre än tjockleken på ett cigarettpapper , i alla fall mellan ordförandeskapets och kommissionens ståndpunkter .
Och det tror jag är allvarligt , framför allt med tanke på rådets kraftfulla ställningstaganden i fråga om Österrike .
Min uppfattning är följande : när det gäller Kina har den förment konstruktiva dialogen inte gett någonting - eftersom vi vet att Europeiska unionens Kinapolitik har misslyckats totalt - men värre ändå är att denna dialog har gett kineserna nya argument för att öka förtrycket , att i än högre grad undertrycka religion och frihet ( vilket Wallström har framhållit på Internet ) , och det i alla områden , i Tibet , det inre Mongoliet och Östturkestan .
Det finns inte ett enda område inom det kinesiska civila samhället där vi inte kan bevittna en tillbakagång .
Detta är ett säkert faktum : Kina är det stora hotet , vårt stora hot , det hot vi måste konfronteras med , ett hot mot freden .
Det är demokratins antites , och ni vet likaväl som jag att kineserna , det kinesiska ledarskapet , är kommunistiskt i första hand och kinesiskt i andra .
Kina älskar att tala med kluven tunga .
Så länge vi inte har en bestämd ståndpunkt kommer vi inte att utverka någonting från de kinesiska myndigheternas sida .
Jag anser därför att vi bör gripa tillfället i flykten .
Vi måste ansluta oss till det amerikanska initiativet .
Vi måste lägga fram en hård text .
Denna text måste röstas igenom .
Vi måste arbeta .
Det krävs att de femton EU-medlemmarna redan i dag arbetar tillsammans med Förenta nationernas medlemsländer , för att ett beslutsamt fördömande äntligen skall uttalas , och för att det sedan , på dessa grunder , skall kunna skapas ett utrymme för dialog .
Herr talman !
Jag skulle vilja försöka anlägga ett annorlunda perspektiv på detta ämne .
Som ni känner till gick i måndags en obemannad luftfarkost in i omloppsbana runt en jordnötsformad asteroid med namnet Eros , som inte är särskilt avlägsen från jorden .
Fotografier visar oss att det inte finns något liv på asteroiden , men mycket längre ut i vår galax , Vintergatan , finns det omkring 300 miljarder stjärnor , många med planeter .
Bortanför Vintergatan finns det omkring 300 miljarder andra galaxer , med oräkneliga stjärnor och planeter .
Det är därför troligt att det finns mängder av liv där ute , som är mycket mer avancerat än vad vi är .
Med tanke på att de första televisionsprogrammen från jorden nu befinner sig 50 ljusår ut i rymden , långt bortom de närmaste stjärnorna , ber jag er att tillsammans med mig föreställa er vad livet där ute tänker om oss när de betraktar oss .
Vad ser de ?
De ser en vacker planet som sprudlar av liv , men de ser dess atmosfär förorenas och värmas upp .
De ser dess skogar huggas ned och öknar spridas ut sig .
Av varelserna kan de se många djur som behandlas grymt , ovanliga arter som utrotas för alltid .
Hur ser de på den just nu dominerande arten - det vill säga på oss ?
Ja , de ser planetens resurser vara ojämnt fördelade .
De ser krig över landområden , medicin mot sjukdomar , men inte i de delar av världen där den bäst behövs , skolböcker - men inte överhuvudtaget i de minst utvecklade områdena av vår värld , 50 procent av världens befolkning ringer aldrig ett telefonsamtal under hela sitt liv .
Vad ser de när de betraktar förhållandet mellan människorna ?
De ser oss döda varandra .
De ser oss begränsa varandras friheter .
De ser en oändlig rad av lokala krig .
De ser några av våra barn värvas till armén som soldater eller utnyttjas som prostituerade eller som slavar .
De ser en ojämlik behandling av män och kvinnor , av människor av olika ålder , av minoriteter , av människor med olika hudfärg , av raser , av religionsanhängare , av invandrare , till och med av grannar .
Vi känner alla till bilden .
FN : s konvention om mänskliga rättigheter för 50 år sedan var ett försök att rätta till detta .
Vi bör hedra det - och jag tycker att vi gör det .
Det är bara i Europa som de mänskliga rättigheterna är lagligt bindande .
Det finns här i Europaparlamentet vissa ledamöter som inte vill att stadgan om rättigheter , som diskuteras för närvarande , skall bli lagligt bindande .
Jag säger : Fy skäms på er !
De mänskliga rättigheterna borde vara lagligt bindande i alla världens länder .
Det är det målet som vi måste arbeta mot .
Mycket återstår , som kommissionär Patten sade , att göra .
Avslutningsvis , om ni frågade mig : Tänk om det inte finns något liv där ute bland stjärnorna , tänk om vi är ensamma ? - vilket är en lika respektingivande tanke - , skulle jag svara : Tycker ni inte att vi har ett ansvar att lära våra barn att uppföra sig väl , innan vi låter dem ge sig i väg för att befolka andra planeter ?
Herr talman !
Mänskliga rättigheter är universella , okränkbara , inbördes beroende och sammanflätade .
Denna berömda slogan , hämtad från slutsatserna från FN : s världskonferens om de mänskliga rättigheterna 1993 kan många utantill .
Det är fint .
Men hur ligger det till med människorättspolitiken inom EU självt ?
Återspeglas denna syn på beroende där ?
Har Europeiska unionen egentligen en människorättspolitik ?
Med denna fråga syftar jag inte på den möda medlemsstaterna har med att samordna sina ståndpunkter i fråga om utrikespolitiken och visa upp en enig linje gentemot kränkningar av de mänskliga rättigheterna på annat håll , exempelvis i Kina .
Nej , herr talman , jag åsyftar avsaknaden av en människorättspolitik inom Europeiska unionen .
I Österrike har en ny regering kommit till stånd där ett politiskt parti deltar som alltid har förkunnat ett budskap som kännetecknas av rasism och intolerans mot minoriteter .
Här hotar således en fara för de mänskliga rättigheter som EU hyllar som en av sina principer , men reaktionerna på dessa händelser har tydliggjort att det saknas en sammanhängande ram inom vilken en lämplig reaktion kan formuleras .
Den allmänt citerade artikel 7 i fördraget , som möjliggör att en medlemsstat där allvarliga och upprepade kränkningar av de mänskliga rättigheterna konstateras kan fråntas sina medlemskapsrättigheter , är naturligtvis bara en sista utväg , det slutliga botemedlet , vilket i fallet med Österrike bara citeras i brist på bättre och som varning .
Det finns därför behov av en fullvärdig människorättspolitik för och av Europeiska unionen , en politik för främjande och tillämpning av de mänskliga rättigheterna inom EU självt .
En sådan politik skulle behöva bestå av ett flertal element .
För det första : det måste finnas en normativ ram där det glasklart står beskrivet vilka rättigheter EU vill säkerställa för sina invånare .
Arbetet med att upprätta en sådan stadga har nu påbörjats , men frågan om rättsstatus och den strategiska betydelsen för detta dokument kan vi inte längre skjuta framför oss eller lägga ut på lärda yrkesjurister .
Detta är en politisk fråga som kräver ett snabbt svar från regeringskonferensen och från parlamentet .
För det andra : det måste utvecklas en skala av instrument som möjliggör en flexible respons och som inte försätter oss i den situationen att vi måste välja mellan en sista utväg och ett slag i luften .
Jag tänker i detta sammanhang på systematisk dokumentation och informationsinsamling , professionella övervakningsformer , utveckling av informationsåtgärder , användning av penningflöden för att stödja demokratiska krafter i det berörda landet , en mer kreativ användning av den multilaterala diplomatins medel , som organiserad dialog och fact finding missions och vad mer hör till .
För det tredje : inom de olika EU-institutionerna måste det tydligt fastställas var ansvaret för människorättspolitiken inom Europeiska unionen ligger och vilka uppgifter och befogenheter det för med sig .
Kommissionen och rådet måste var och en för sig redan ut begreppen vad det beträffar .
För parlamentet behövs inte detta längre , med tanke på att det i vår arbetsordning fastställs att utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor har dessa befogenheter .
Men då är det ändå underligt att den resolution som skall avsluta denna debatt om de mänskliga rättigheterna har förberetts i parlamentets utrikesenhet och att det utskott som jag nyss nämnde , och som jag själv utgör en del av , inte har kommit ifråga .
Herr talman !
Parlamentet är rubbat och splittrat .
Med tanke på vår trovärdighet bör vi tala med en röst och inte behöva låtsas som om mänskliga rättigheter inom EU är någonting annat än mänskliga rättigheter på andra håll i värden .
Jag tror att detta också skulle kunna vara till nytta för vår trovärdighet i FN : s kommission för mänskliga rättigheter .
Herr talman !
Vad krävs det för att diskussionen om de mänskliga rättigheterna skall bli någonting annat än vad den är i dag : ett ideologiskt instrument som medverkar till folkens träldom och inte till människors frihet ?
Vi måste först och främst gå tillbaka - bortom människan själv , som inte är universums härskare - till källan för all verklig rätt och civilisationens grundläggande värden , förutan vilka de eviga kraven på rättigheter alltid slutar i tyranni , i blodigt tyranni .
Med hela den europeiska antika och medeltida traditionen måste vi gå tillbaka till universums naturliga ordning , dvs. skapelsen , och antagligen bortom den , till skaparens planer .
Då skulle vi bli varse att barnets rättigheter endast respekteras inom en riktig familj , att arbetarens rättigheter endast respekteras inom ekonomins mellanled , som man nyss har förstört , och att medborgarens rättigheter endast respekteras inom suveräna nationer .
För det andra krävs det att doktrinen om de mänskliga rättigheterna inte längre instrumentaliseras , på det sätt som sker i dag , till en ideologisk krigsmaskin i händerna på en exklusiv elit som tillskansar sig rätten att ensidigt förordna om vem som företräder de mänskliga rättigheterna och vem som står utanför deras sfär , vilket gör att de kan förneka all legitimitet och , vid behov , all frihet för dem som den likriktade tanken har pekat ut som politiskt inkorrekta .
Ingen frihet för frihetens fiender , det sade företrädarna för det revolutionära skräckväldet för 200 år sedan , den revolution som tyvärr blev en förebild för alla moderna former av totalitarism .
Inga mänskliga rättigheter för de mänskliga rättigheternas fiender , det säger i dag de som lovprisar den nya världsordningen , de som nästan helt och hållet regerar finansiella sammanslutningar , internationella institutioner , nätverk på medie- och kulturområdet , pedagogiska institutioner och jag vet inte allt .
Vad återstår till exempel av österrikarens rätt att fritt välja sitt öde , om hans val dikteras av dem som i hans ställe beslutar om vad som är passande eller inte passande att göra , och om hans ledare - valda genom en legal och legitim process - tas emot på ett förolämpande sätt , som när de nyligen togs emot av er , herr rådsordförande , herr minister från Portugal .
Jag vet inte om han är här för att lyssna på mig .
Vad återstår det av de mänskliga rättigheterna för dem som sympatiserar med partiet Vlaamsblok , ett av de största partierna i den flamländska regionen , om det belgiska parlamentet i morgon antar det osannolika , ovärdiga och vanhedrande lagförslag som kommer från dess huvudsakliga politiska konkurrent , partiet Volksunie , ett förslag som endast syftar till att tillintetgöra rivalen ?
Vad återstår av rätten till en kritisk granskning av vår historia , när författare och utgivare förföljs , vilket hände så sent som i går i appellationsdomstolen i min stad Lyon , då den unge historikern Jean Plantin utsattes för absurda , arroganta och kränkande anklagelser från generaladvokaten Jean-Olivier Viout , ett belåtet uttryck för den likriktade tanken och intellektuell konformism ?
Vilken märklig uppfattning om de mänskliga rättigheterna är inte detta : att svekfullt förväxla fredlig patriotism med krigisk nationalism ; legitima protester mot invandringspolitiken med jag vet inte vilken typ av främlingsfientlighet , och det nödvändiga försvaret av identiteter med rasism !
Vilka mänskliga rättigheter har de miljoner fransmän som röstar på Nationella fronten , människor som har berövats alla sina politiska företrädare och som dagligen svärtas ned , till exempel i måndags i den statstelevision som de tvingas betala för via skattsedeln , då ett rättframt men med rätta förbittrat uttalande av en av våra kolleger , Le Pen , får tjäna som förevändning för orättfärdiga fördömanden - vilket utgör ett brott mot lagen , ett brott mot rättvisan , rättrådigheten och moralen - och då man i dag , i strid med de allra tydligaste föreskrifter , gör anspråk på att beröva denne företrädare det mandat han har erhållit genom miljoner medborgares röster , och inte genom maktens favör .
Kort sagt , mina kära kolleger , jag kommer att tro på era tal om de mänskliga rättigheterna i Europa när ni tillerkänner era politiska motståndare samma rättigheter som ni beviljar er själva .
Jag kommer att tro på ert tal om de mänskliga rättigheterna i Kina när ni pekar ut den verkliga orsaken till det onda , dvs. kommunismen .
Lyssna till Solsjenitsyns mäktiga röst i hans brev till amerikanerna ; den främsta orsaken till västländernas svaghet ligger enligt honom i en sjukligt uppförstorad lagstadgad individualism , en individualism som långtifrån tillåter enskilda människor att utvecklas , utan i stället banar vägen för en kommande diktatur .
Och det kommer att bli den värsta av diktaturer , eftersom de förslavade inte ens kommer att vara medvetna om sin fasansfulla träldom .
Herr talman !
Principen om de universella mänskliga rättigheterna är otvivelaktigt ett av de viktigaste politiska arven från 1900-talet .
Förintelsen gav för femtio år sedan anledning till att fastställa ett antal grundläggande rättigheter och friheter .
Sedan det kalla kriget upphört har efterlevnad av de mänskliga rättigheterna också blivit ett villkor för internationellt samarbete .
Ledare som kränker dessa principer konfronteras nu med internationell kritik , sanktioner eller till och med rättegång som före detta diktatorer som Pinochet har fått erfara .
Denna utveckling är hoppingivande .
Men den hindrar inte att tillståndet för de mänskliga rättigheterna i världen fortfarande är mycket oroande .
Det är framför allt i krigssituationer som civila skonas allt mindre .
Det förefaller motsägelsefullt .
Aldrig tidigare i historien har den humanitära rätten varit så väl utbyggd .
Aldrig tidigare har så många internationella fördrag varit ratificerade av så många länder .
Ändå förekommer förbrytelser mot de allra mest grundläggande uppförandekoderna i stor omfattning , och det krävs fler civila offer än för ett århundrade sedan .
Kvinnor våldtas systematiskt .
Barn tvångsrekryteras och sätts in i striden .
Övergrepp är inte längre undantag ; de har tyvärr blivit regel .
Det gäller i dag för inte mindre än trettio konflikter över hela världen .
För sen , för selektiv och för splittrad , så skulle man kunna beskriva världssamfundets människorättspolitik .
För sen .
Såväl i Rwanda som i Kosovo visade det sig att FN , trots de många varningarna , kom sättandes för sent och blev en maktlös åskådare till massakrerna , vilket president Havel sagt här under eftermiddagen .
Men inte heller femtio år senare lyckas vi att förhindra folkmord .
Det är således högst angeläget att ägna mer uppmärksamhet åt övervakning och konfliktförebyggande .
Uppsikt över vapenhandeln och en bättre kontroll av medierna är väsentligt i detta ärende .
Människorättspolitiken är också för selektiv .
Natos bombningar av Kosovo under flera månader och medlingsförsöken i Mellanöstern står i bjärt kontrast till den internationella likgiltigheten i fråga om konflikterna i Afrika .
Jag kan inte bli kvitt intrycket av att när det handlar om mänskliga rättigheter , då står inte Afrika högst upp på det portugisiska ordförandeskapets dagordning trots all retorik .
Det är något som jag verkligen beklagar .
Det är inte utan anledning som afrikanerna får intryck av att de är mindervärdiga världsmedborgare .
Jag skulle vilja varna för en försvagning av normerna vid bedömningen av situationen för de mänskliga rättigheterna i Afrika , varvid man börjar betrakta kränkningarna där som något oundvikligt .
Men människorättspolitiken är framför allt för splittrad .
Vi lyckas inte att fastställa en gemensam strategi inom de internationella gemenskaperna , och inte ens inom Europa .
Ta nu Sudan .
Världssamfundet sänder ut motstridiga signaler till det landet .
England öppnar åter sin ambassad i Khartum .
Kanada bjuder in sudaneserna till fredssamtal .
Europa sätter rebellerna i söder under tryck för att få förhandlingar till stånd , och samtidigt börjar amerikanerna isolera regimen och stödja rebellerna militärt .
Det behövs mer samordning , mer informationsutbyte och ett mer samstämmigt handlande där man undviker varje överbud .
Det är bara på det sättet som vi kan följa grundläggarna av den allmänna förklaringen om mänskliga rättigheter på ett konsekvent sätt .
Herr talman !
Jag skulle vilja börja med att säga att om ord kunde lösa problemen , skulle vi alla kunna packa ihop och åka hem .
Men samtidigt som vi i dag talar inne i denna kammares säkerhet , äger tyvärr kränkningar av de mänskliga rättigheterna rum runt om i den fria världen .
Ibland hör vi mindre ju mer vi talar - motioner : ord ; konventioner : ord ; fördrag : ord - , och om vi inte är försiktiga , blir orden själva ett substitut för verklig handling .
Ord inramade i allomfattande och utförliga dokument blir fördrag och konventioner som ofta visas upp som bevis på att ett land respekterar och håller sig till de mänskliga rättigheterna .
Men talade , skrivna eller undertecknade ord är inte i sig själva tillräckligt .
Se på undertecknarna av konventionerna om mänskliga rättigheter och minoriteter , och jämför därefter hur sådana minoriteter , grupper och individer behandlas - listan är skamlig och generande .
Finns det någon som med den minsta trovärdighet kan hävda att kvinnor behandlas jämlikt och rättvist , att barn har mänskliga rättigheter eller att människor inte diskrimineras på grund av sin religion , sin tro , sitt kön , sitt handikapp , sin ålder , sin sexuella läggning , sina åsikter , sin politiska tillhörighet osv . ?
Förtalet av minoriteter i dagstidningar och i andra medier ger bränsle åt diskrimineringen .
Även inom EU utsätts medborgarna fortfarande för kränkningar av de mänskliga rättigheterna och brott mot våra konventioner .
I pressen används dagligen felaktig information och oriktiga framställningar för att förvägra minoriteter jämlikhet inför lagen och för att svärta ned etniska minoriteter .
Uppriktigt sagt har en förtryckarhierarki skapats .
Och så länge som människor inte är jämlika inför lagen , kommer denna ojämlikhet att leda till diskriminering , och de mänskliga rättigheterna kommer att undergrävas .
I vår utvidgningsprocess har vi i EU med rätta lagt tonvikten på mänskliga rättigheter och skydd av minoriteter .
Vi får inte göra avkall på detta åtagande .
Men vi måste också hålla upp spegeln framför oss själva och erkänna våra egna brister .
Ja , konventioner har undertecknats , men det behövs handling .
Jag skulle föreslå er en fortgående granskning av hur de mänskliga rättigheterna tillämpas , en ständig övervakning , inte bara utanför våra gränser , utan också innanför .
Det är av den anledningen som jag skulle välkomna en årlig medlemsstatsrapport från varje enskild stat , i vilken alla anklagelser mot staten liksom de vidtagna åtgärderna skulle tas upp .
För vad som händer i varje medlemsstat händer var och en av oss .
Vad som händer i en annan del av världen påverkar oss .
Pinochet i Chile är lika relevant som Haider i Österrike .
Mänskliga rättigheter och medborgerliga friheter är oupplösligt sammanlänkade .
Mänskliga rättigheter existerar inte isolerat , de hänger samman med vår utvecklingspolitik , vår ekonomiska politik , vår inrikespolitik , de är i själva verket i centrum av våra demokratiska funktioner .
Jag skulle vilja upprepa vad Patten sade : Vi måste engagera oss , vi måste informera och utbilda och därigenom få till stånd en verklig och bestående förändring .
Herr talman ! "
Europa står för ideal , värderingar och principer .
Vi måste lyfta fram Europas andliga historia .
Gemensamt måste vi återupprätta de värderingar som enar Europa .
Andliga värden har spritts från Europa ut över hela världen .
Vi måste leva med våra samveten . "
Så sade för tre timmar sedan Tjeckiens president Vaclav Havel i denna kammare .
I ett synnerligen upplyftande tal , präglat av människokännedom , vishet , historisk kunskap och insikt om Europas andliga och kristna arv , pekade han på inspirationskällor för vårt arbete kring människans värde och kring människorätten .
Vi skall vara tacksamma för att det finns statschefer som Vaclav Havel i vårt Europa .
Jag vill ta upp två saker .
Det gäller först det civila samhället .
Vaclav Havel nämnde att i Östeuropa slog kommunistregimerna metodiskt sönder det civila samhället : folkrörelserna , kyrkorna och de oberoende fackföreningarna .
Detta sker i Kina med Falun Gong-rörelsen och med de katolska och protestantiska kyrkorna .
Det sker med lamaismen i Tibet .
Vi får aldrig glömma bort försvaret av det civila samhället .
Jag vill också ta upp dödsstraffet .
EU , liksom mitt land Sverige , bygger sin människosyn på det lika , unika och okränkbara människovärdet .
Utifrån denna princip skall människan alltid ha en chans att komma tillbaka .
Säg det till Förenta staternas regering , till Rysslands regering och till Kinas regering !
Herr talman !
Herr rådsordförande !
Herr kommissionär !
Jag anser att EU-medlemsstaternas strategi i Genève bör vara att prioritera situationen i Kosovo , Mexiko , Saudiarabien , Sierra Leone och Kina .
Vad Kina beträffar bör vi inte låta bli att ta upp frågan bara för att diskussionen om den kan bli blockerad .
Det är dock av högsta vikt att EU talar och agerar som en enhet , och hot om handelssanktioner bör snarare stärka än försvaga vår beslutsamhet .
Om de beslut som slutligen kommer att fattas i Genève skall ges sitt fulla uttryck , måste den höga kommissionären för mänskliga rättigheters kontor emellertid förses med de nödvändiga resurserna .
Förenta nationernas ekonomiska resurser är utspridda i ett mycket tunt lager , och många centrala program är därför beroende av frivilliga bidrag för att kunna fungera .
Resurser behövs också för att främja praktiskt samarbete och mänskliga rättigheter , för strategisk planering , för att fastställa prioriteringar och för att stärka kommunikationen mellan givarsamfundet och Förenta nationernas medlemsstater .
Därför framförde nyligen den höga kommissionären en vädjan om 53 miljoner US-dollar årligen för att göra det möjligt för sitt kontor att utföra dessa uppgifter .
Europeiska unionen och dess medlemsstater bör ta täten och tillhandahålla en betydande andel av dessa medel .
Genom att göra det skulle vi inte bara genera Förenta staterna och därigenom få landet att axla sitt ansvar i fråga om FN-finansieringen , utan vi skulle också bevisa att våra utfästelser om att försvara de mänskliga rättigheterna är mer än bara tom retorik .
Herr talman !
I denna debatt handlar det framför allt om förberedelserna inför FN : s årliga session om de mänskliga rättigheterna inom kort och om kommissionens och rådets insatser i det sammanhanget .
Låt mig först och främst säga att jag är mycket nöjd med det som har tagits upp hittills av Patten och av ministern , och jag tycker också att det är positivt att såväl Kina som Kuba tas upp till diskussion .
Kuba är fortfarande den sista diktaturen i Sydamerika , och det får vi inte glömma bort med tanke på all sympati för Kuba som här och där gör sig gällande .
Det är en diktatur och således ingen demokrati .
Jag vill under mina två minuter be om uppmärksamhet för två länder som jag har ett särskilt band till .
Det är i första hand Indonesien .
Vi är naturligtvis mycket glada över att Indonesien har en ny regering och att Wahid och Soekarnopoetri innehar posterna som president och vicepresident .
Vi gläder oss också åt att situationen i Timor sakta men säkert går i rätt riktning .
Men jag vill tala om för er att på Moluckerna , ett område som ligger alldeles ovanför Timor , är våldet fortfarande inte under kontroll .
Där har tusentals dödsoffer krävts under de senaste två åren .
Tiotusentals människor är på flykt .
Man har inte fullständig kontroll över händelserna .
Jag vet att det i morgon eller i övermorgon kommer ett stort program på nederländsk TV där man vädjar om observatörer , bara för att observera precis det som sker där så att det som har skett i varje fall blir registrerat , även för framtiden , för människorättskommissionerna .
Min angelägna vädjan är , och det är också en punkt som ett flertal gånger har fastlagts här i resolutioner : kan ni inte förhandla så att observatörer skickas till Moluckerna ?
Tusentals döda , tusentals sårade , tiotusentals på flykt borde väl vara tillräckligt .
Mitt andra land , och där kommer jag att fatta mig mycket kort , för Patten känner till det mycket väl , är Burma .
Det kan ändå inte gå för sig att vi tiger om Burma .
Jag har en känsla av att det landet sakta men säkert faller i glömska .
Sedan tio år tillbaka finns där en vald president som sitter i husarrest .
Sedan tio år tillbaka fungerar inte parlamentet längre .
Otaliga parlamentsledamöter har dödats eller flytt , och det är bara några enstaka som bor kvar i Burma .
Det finns hundratusentals flyktingar från Burma i Thailand och Indien , och ändå verkar det som om landet inte längre får någon uppmärksamhet .
Jag anser , i synnerhet i förlängningen av vändningen i Indonesien , att även Burma återigen måste sättas upp på dagordningen .
Det går ju inte för sig att Aung San Sui Kyi känner sig helt lämnad i sticket , även av Europa .
Min vädjan är egentligen att även det landet på nytt skall sättas högt upp på dagordningen .
Herr talman , herr tjänstgörande rådsordförande , ärade kommissionär !
Europeiska unionens roll i världen får inte avgöras enbart genom ekonomisk makt .
Det är viktigt att vi också utmärker oss när det gäller kampen för de mänskliga rättigheterna , vare sig det gäller från vår sida eller dem som vi står i förbindelse med .
Europaparlamentet har stått i centrum för kampen för de mänskliga rättigheterna , man har lyckats se bortom egoism och " nationella intressen " som många gånger har orsakat motsättningar länderna emellan och till och med mellan Europeiska unionens institutioner .
Man kan exempelvis konstatera att Europaparlamentet aldrig glömde situationen i Östtimor , något som hade varit fatalt för en rättvis lösning för folket , ett folk som alltid motsatte sig den indonesiska ockupationen .
Det var inte länge sedan som vi därför motsatte oss försäljningen av vapen till Indonesien , en ståndpunkt som rådet tyvärr inte tog i beaktande .
Det är inte tillräckligt att bara försöka hindra upprörande aggressioner av människor eller institutioner mot de svaga .
De gärningsmän som begått kränkningarna får under inga omständigheter gå ostraffade , oavsett vem det är och var det är , i Indonesien eller i Angola , i Kuba , i Kina eller i Burma , och oavsett om gärningsmannen är en civilperson eller en militär , en general eller en minister .
Rättvisa måste skipas i Indonesien .
Rättvisa måste skipas i Östtimor .
President Wahid behöver vårt stöd för att klara av den svåra situation han befinner sig i .
Efter påtryckningar av PPE tog man i sista minuten uttryckligen med Östtimor i resolutionen .
För det som hände där , och som jag som företrädare för Europaparlamentet delvis fick tillfälle att se , måste någon ställas till svars och bestraffas .
När vi talar om Östtimor måste vi också komma ihåg situationen med tiotusentals flyktingar från Östtimor på indonesiskt territorium , i en omänsklig situation , kontrollerade av indonesisk militär och milis och använda som påtryckningsmedel .
Det är en outhärdlig situation som vi snabbt måste sätta stopp för .
Herr talman !
I egenskap av rådets ordförande vill jag i all korthet påpeka att ordförandeskapets arbete framför allt går ut på samordning , att försöka nå en gemensam ståndpunkt för de initiativ som de femton måste anta i rådet .
Erfarenheter från tidigare sessioner i utskottet för mänskliga rättigheter har visat - just på grund av ordförandeskapens samordningsförmåga - att Europeiska unionen har lyckats stärka sin roll som organisation med egen politik i kommissionen , vilket är det viktiga .
Jag vill också säga att Europaparlamentets delaktighet i de förberedande arbetet är viktigt för en samordnad bekräftelse av Europeiska unionens ståndpunkter .
Ordförandeskapet tar därför givetvis gärna emot alla förslag och bidrag till de två resolutioner som har lagts fram här .
Jag vill också påpeka att många av ledamöterna menade att de mänskliga rättigheterna skall vara en central del i den europeiska identiteten och att respekten för de mänskliga rättigheterna skall ses som en grundläggande princip för det internationella samarbetet från Europeiska unionens sida .
Därför måste vi samordna den europeiska politiken om mänskliga rättigheter på ett bättre sätt , vilket gör att vi måste klargöra våra ståndpunkter och klart och tydligt tala om vilka situationer som vi anser vara de mest oacceptabla , till exempel den i Kina som många av ledamöterna refererade till .
Vi kunde också notera den oro andra ledamöter känner inför situationer i andra länder , må vara i Indonesien eller i Timor , i Moluckerna eller i Burma .
Avslutningsvis vill jag särskilt kommentera ledamot Van Heckes anförande om de mänskliga rättigheterna i Afrika och portugisiska ordförandeskapets roll och prioriteringar , där han ifrågasätter vår uppriktighet när det gäller hur det portugisiska ordförandeskapet prioriterar relationerna med Europeiska unionen .
Jag vill bara säga att det portugisiska ordförandeskapet under dessa två månader för första gången har kunnat genomföra ett ministerrådsmöte ( utvecklingssamarbete ) vars agenda , må vara informellt , dominerades av förbindelserna Europeiska unionen-Afrika - och att det var detta som fick de femton ministrarna att sammanträda i Lissabon för att debattera den nya dimensionen av de nya förbindelserna - och jag kan inte låta bli att påpeka att vi faktiskt har avslutat de viktiga förhandlingarna om den nya konvention som skall ersätta Lomékonventionen , och att vi trots svåra förhandlingar har lyckats förbereda genomförandet av det första toppmötet Europeiska unionen-Afrika .
Det var anledningen till att jag inte kunde låta bli att besvara ledamot Van Heckes fråga . .
( EN ) Herr talman !
Det har varit en mycket nyttig debatt .
I ett eller två tal har särskilda frågor som vi gör klokt i att överväga mycket noga tagits upp .
Till exempel tog Maij-Weggen upp både Indonesien och Burma , och hon sade några viktiga saker om dessa båda länder och om situationen för de mänskliga rättigheterna där .
Vad jag skulle vilja koncentrera mig på helt kort är en eller två röda trådar som har löpt genom vår debatt .
En av de allra första talarna , Wuori , talade om de kommentarer som Havel gjorde tidigare i dag .
Det var ett anmärkningsvärt tal , och jag hoppas att även Gollnisch , som inte har möjlighet att vara med oss nu , kunde höra detta tal .
Jag hoppas också att , om det finns något liv i yttre rymden , vilket Newton Dunn spekulerade i , även dessa varelser fångade in Havels tal .
Havel påminde oss om att unionen inte bara handlar om marknader , om BNI-tillväxt , utan att det är en union av värderingar , som avspeglas i fördragen och som avspeglas i våra åtaganden på hela området för externt bistånd , som avspeglas ganska tydligt i de uppgifter som vi har fått i uppgift att utföra .
Hur genomför vi det som föreskrivs i fördragen i alla dessa ord om utvecklingsbiståndsprogram ?
En eller två ärade medlemmar , Ferber och Cushnahan , talade om gapet mellan retorik och verklighet .
Cashman sade , vilket på sätt och vis är riktigt , att ord inte är ett substitut för verklig handling .
Ord kan , naturligtvis , ge en viss effekt , vilket Malmström gav exempel på .
Hon sade att hon har mottagit ett brev från Kinas ambassadör , en mycket älskvärd och intelligent man som företräder och arbetar för sitt land , i vilket han talar om att hon har fel och att Europaparlamentet har fel i sin syn på de mänskliga rättigheterna i Kina .
Jag tror att hon efter sitt tal kommer att få ta emot en störtflod av brev från de kinesiska myndigheterna .
Hon kommer att kunna fylla ett dokumentskåp med brev om vad som hävdas vara den verkliga situationen i Kina .
Jag tror att hon återgav åsikterna hos många icke-statliga organisationer , hos många människor som beundrar den kinesiska civilisationen men som är bekymrade över vad som händer i Kina i dag .
Det är naturligtvis helt rätt av vi måste överväga handlingar , och i det allra första talet av Salafranca nämndes två saker , bortsett från Genèvemötet , som utgör handlingar , av vilka en naturligtvis möjliggörs av Europaparlamentets , på de europeiska skattebetalarnas vägnar , generositet - det vill säga den budget som vi kan använda på verksamhet som hör samman med de mänskliga rättigheterna , omkring 100 miljoner euro som används genom program , för vilka jag är ansvarig , och som huvudsakligen går till icke-statliga organisationer för att främja mänskliga rättigheter och demokratisering .
Vi kommer med parlamentet att vilja dela , som vikarierna säger , våra åsikter om hur detta utgiftsprogram för att stödja mänskliga rättigheter bäst kan fokuseras och bäst kan riktas in under de kommande åren .
Dessutom har vi den fråga som togs upp av Salafranca , som jag beklagar inte kan vara här med oss i slutet av denna korta med nyttiga debatt .
Dessutom har vi frågan om vår övergripande politik om mänskliga rättigheter och förhållandet mellan de mänskliga rättigheterna och utrikespolitiken .
Jag vill påminna parlamentet om att kommissionen före halvårsskiftet kommer att offentliggöra ett omfattande intellektuellt förslag om att placera de mänskliga rättigheterna i hjärtat av den gemensamma utrikes- och säkerhetspolitikens utveckling .
Det är oerhört viktigt , och om jag inte redan hade tyckt det , skulle jag efter att ha lyssnat till Havels anmärkningsvärda tal tidigare i dag utan tvekan ha kommit fram till den slutsatsen .
Det har varit en nyttig debatt .
Jag hoppas att vi kan ha flera debatter som denna .
Jag hoppas särskilt att vi kan ha debatter om några av de sätt på vilka vi kan omsätta dessa goda föresatser i praktisk handling på de platser där det behövs , där människor ännu torteras , där människor ännu våldtas och ännu nekas den slags medborgerliga rättigheter som denna kammare - liksom jag - tar för givna .
Jag har till följd av detta uttalande fått 7 resolutionsförslag i enlighet med artikel 37.2 i arbetsordningen .
Härmed förklarar jag debatten avslutad .
Omröstningen kommer att äga rum på torsdag .
 
Cypern och Malta Nästa punkt på föredragningslistan är debatten om : rådets uttalande om Europeiska unionens inställning till utvecklingen av Cypernfrågan ; betänkande ( A4-0029 / 2000 ) av Brok för utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik om förslaget till rådets förordning om genomförande av åtgärder inom ramen för en strategi inför anslutningen till Cypern och Malta ( KOM ( 1999 ) 535 - C5-0308 / 1999 - 1999 / 0199 ( CNS ) ) .
Jag överlämnar ordet till Seixas da Costa , som företrädare för rådet .
Herr talman , ärade kollegor !
I egenskap av Europeiska unionens rådsordförande vill jag informera om de återupptagna cypriotiska förhandlingarna och vad som där skett .
Jag tror att det är uppenbart för oss alla att det som hände i Helsingfors i slutet av förra året och den nya stämningen i förbindelserna mellan Europeiska unionen och Turkiet återspeglar en grundval på gemenskapsplanet som inte kan låta bli att påverkas av förbindelserna mellan de två samfunden på Cypern .
Jag vill också framhålla att i fjol , i början av december , ägde den första förhandlingsrundan rum i New York , förhandlingar som under många år varit avbrutna mellan de båda cypriotiska samfunden på norra och södra delen av ön .
De samtal som fördes var av indirekt natur med medlaren Álvaro de Souto som Förenta nationernas särskilda sändebud .
Nya förhandlingar ägde rum i januari i år , från och med den 31 januari , och en tredje runda beräknas börja den 23 maj i New York .
Möjligheten finns , även om detta på intet vis har bekräftats , att samtalen kan fortgå direkt och fortlöpande fram till september i år .
Det väsentliga i den här diskussionen kan sammanfattas i fyra punkter : Säkerhetsaspekten , regeringsstrukturen , territoriella justeringar samt flykting- och skadeståndsfrågorna som härrör från den situation som uppstod efter öns delning .
Man hade kommit överens om att inkludera andra frågor och därför har företrädaren från öns norra del , Rauf Denktash , föreslagit följande : frågan om suveränitet , förtroendeskapande åtgärder samt frågan om att lyfta embargot på de produkter som kommer från norra delen .
Av de samtal som hittills har förts har i huvudsak följande uppnåtts : man skissar på möjligheten att skapa en direkt informationskanal mellan Europeiska unionen och öns norra del , utan att detta nödvändigtvis betyder att man på det internationella planet erkänner den delen av ön som en juridisk person med syfte att underlätta ett antagande av gemenskapsrätten vid en eventuell anslutning av hela ön , om man under tiden har lyckats finna en global lösning på problemet med öns delning .
Det andra som uppnåtts och som vi anser är betydelsefullt är det uttalande som gjordes av Förenta nationernas generalsekreterare i slutet av andra dagens samtal .
Han menade att om man lyckades lösa problemet globalt så skulle en sådan innebära att norra delen av ön erkänns med sina särdrag .
Detta är den ståndpunkt som generalsekreteraren intog och som vi måste beakta i vår framtida analys .
Man har vissa förväntningar på den tredje förhandlingsrundan tack vare de bakgrundsförslag som håller på att förberedas och där företrädare från Förenta staterna och Förenade kungariket deltar , i första hand när det gäller säkerhetsfrågor och den författningsenliga strukturen , frågor som , för det andra , förmodligen kommer att presenteras av Förenta nationernas generalsekreterare under de här samtalen , något som kommer att inträffa efter de val som förrättas i norra delen av ön den 18 april .
Europeiska unionens portugisiska ordförandeskap följde exemplet från tidigare ordförandeskap och beslutade sig för att utse en företrädare för att hålla kontakt med de parter som är involverade i frågan .
Företrädaren har redan kontaktat parterna och har i nära samarbete med Förenta nationernas generalsekreterare följt arbetet under de olika förhandlingsrundorna .
Det är i första hand vår avsikt att fortsätta profilera Europeiska unionen i den här frågan , i synnerhet när man kan konstatera att Cypern vill ansluta sig till Europeiska unionen medelst ett ganska framfusigt förhandlingsförfarande , något som givetvis väcker förhoppningar och samtidigt avgör om Europeiska unionen skall ha någon roll av betydelse i det här sammanhanget .
Diskussionens inriktning och vårt deltagande i samma diskussion har i huvudsak bestått i att utnyttja ett något lugnare klimat skapat av övertygelsen , något som vi alla delar , att det är nödvändigt att fortsätta förhandla och att fortsatta förhandlingar och bevarad rytm i sig är avgörande för förhoppningen om en slutlig lösning .
Det finns en annan fråga av vikt , jag refererade till den i början av mitt uttalande , som har att göra med Turkiets iver att bidra till förberedelserna för en anslutning av norra delen av ön .
Vi menar att vi inte bara måste läsa Europeiska rådets slutsatser från Helsingfors med viss noggrannhet utan också med försiktighet , samtidigt som vi måste följa det som kan vara de turkiska myndigheternas tillgänglighet för att bidra till att lösa den här frågan .
Jag var själv i Ankara där jag fick tillfälle att tala med premiärminister Bülent Ecevit om detta , och trots det faktum att vi är medvetna om såväl svårigheterna som särdragen och turkarnas överdrivna känslighet i den här frågan , så anser jag att en möjligheternas dörr har öppnats som måste tas tillvara .
Denna möjligheternas dörr behöver en kombination av faktorer , en av dem , och det är ingen mening att dölja det , har att göra med själva dynamiken i förbindelserna mellan Turkiet och Europeiska unionen .
Grundläggande för den här frågans framtid .
Å andra sidan menar vi att det är viktigt att informationsutbytet mellan kommissionen och cyprioterna i norr uppmuntras , utan att , och låt detta klargöras , utan att detta medför något som helst formellt erkännande , vilket fortfarande har att göra med hur Europeiska unionen ställer sig i den här frågan Vi menar dock , och jag tror att även kommissionen har tolkat det så , att hela förfarandet med ett närmande till gemenskapsrätten i riktning mot ett globalt integrationsförfarande av ön inom ramen för Europeiska unionen vid en framtida anslutning , innebär att norra delen av ön , så snart som möjligt , måste involveras samtidigt som Europeiska unionen också måste få tillgång till den information som kan ge substans åt själva anslutningsprojektet i sina bemödanden att utvärdera villkoren för en anslutning .
Å andra sidan innebär det att vi från rådets sida måste se till att kommissionen engagerar sig , vilket också parlamentet kan göra .
Jag tror att vi måste visa kommissionen vårt förtroende när det gäller den roll man skall spela .
Å andra sidan : med hänsyn till hur skickligt , intelligent och kompetent generalsekreteraren har drivit de här förhandlingarna och försökt bidra till en harmonisering av parternas ståndpunkter samt med hänsyn till Förenta nationernas inre struktur så tror jag slutligen , precis som ordförandeskapet , att vi aktivt måste fortsätta att samarbeta med Förenta nationerna .
Som jag inledningsvis sade så kan man konstatera att slutsatserna från det europeiska toppmötet i Helsingfors i december förra året fick ett stort inflytande på utvecklingen av parternas ståndpunkter i förfarandet .
Regeringen i Nicosia sade sig vara nöjd med slutsatserna från Helsingfors , vilka öppnar dörren till en anslutning till Europeiska unionen utan att på förhand ha löst öns delning .
Jag kan emellertid inte låta bli att notera att samma myndigheter är oroade över eventuella påtryckningar för att lösa de frågor som uppstår i och med en delning , frågor som uppenbart kommer att innebära en del eftergifter .
Det här har att göra med den utveckling man kunnat notera när det gäller förflyttning av befolkningen och möjligheten att omorganisera en förflyttning av samma befolkning i fall man når en annan överenskommelse för ön .
Å andra sidan är cyprioter och turkar rädda för att Turkiets kandidatur till Europeiska unionen kan komma att leda till ökad medgörlighet från Ankaras sida i den här frågan , något som inte är lönt att dölja .
Oberoende av om det i de båda gemenskaperna finns en tendens till misstro inför ett sådant närmande , så tror jag att de aspekter som kan få myndigheterna på båda sidor att negativt tolka situationen , också kan vara de grundläggande skälen till förhoppningen om en slutgiltig lösning .
En sådan slutgiltig lösning kommer givetvis att färgas av en av de viktigare händelserna på området under den här perioden , nämligen den synnerligen positiva utvecklingen av förbindelserna mellan Aten och Ankara och den utomordentligt viktiga roll utrikesministrarna här spelade , såväl George Papandreou som den turkiske utrikesministern Ismail Cem .
Vi tror att villkoren för en positiv utveckling har skapats .
Från vår sida , från rådets ordförandeskaps sida , kommer vi att fortsätta att uppmärksamma utvecklingen , vi kommer att fortsätta att samarbeta med generalsekreteraren och med dennes personliga sändebud i den här frågan .
Vi kommer att informera gemenskapsinstitutionerna om vad vi kan göra och vad som skulle kunna göras när det gäller samordning , inte bara på det politiska planet utan också vad kommissionen med sina befogenheter kan åstadkomma inför anslutningsförfarandet , och vi kommer särskilt att berätta om den flexibilitet som parterna visade prov på i den här frågan .
Herr talman , ärade damer och herrar !
Debatten i dag befattar sig med en fråga som är särskilt viktig ur två synvinklar .
Först är det fråga om finansieringen för att Cypern och Malta fullt ut skall kunna omfattas av förberedelsestrategin för medlemskap .
Men det handlar även alldeles särskilt om fredsprocessen på Cypern och därmed även om stabilitet och säkerhet i Medelhavsområdet .
Jag vill inleda med att säga några ord om den budgetförordning som kommissionen lade fram för Cypern och Malta i oktober förra året .
Jag är ytterligt tacksam mot Brok , föredraganden och ordföranden i utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik , för dennes betänkande , som bildar en utmärkt grund för våra överläggningar i dag .
Vi behöver detta instrument .
Det ersätter de finansprotokoll som löpte ut i slutet av 1999 .
Vi behöver dessa instrument för att kunna fullgöra våra finansiella förpliktelser när det gäller förberedelsestrategin för Malta och Cypern .
Jag är mycket tacksam över att parlamentet stöder kommissionen i dess strävan att slutbehandla och godkänna förslaget till förordning så snabbt som möjligt .
Utskottet för utrikesfrågor samt budgetutskottet har lämnat in en rad ändringsförslag .
En del av dem kan kommissionen acceptera .
Det finns två punkter som jag gärna vill yttra mig om , två punkter som jag vet ligger parlamentet särskilt varmt om hjärtat .
Det ena gäller finansieringen som sådan : hur mycket pengar skall vi då alltså egentligen satsa ?
Kommissionen kommer att föreslå en finansiering i storleksordningen 95 miljoner euro .
Även rådet har enats om denna siffra .
Jag vet att parlamentet önskar en mer omfattande finansiering , och jag kan också förstå varför .
Tro mig , som ansvarig ledamot av kommissionen skulle även jag gärna ha mer pengar till förfogande för detta ändamål .
Men situationen är nu en gång sådan att man för tillfället inte kan enas om ett högre belopp .
När allt kommer omkring är det ändå budgetmyndigheten som måste fastslå det slutgiltiga beloppet .
Den andra frågan som är av vikt gäller hur de ekonomiska medlen under rubrik 7 i budgeten skall användas .
Detta är ju endast skenbart en teknisk fråga .
I högsta grad är det en politisk fråga .
Jag själv har vid ett annat tillfälle redan sagt att jag anser detta vara en korrekt tanke .
Jag tror mig kunna säga - utan att kommissionen för den skull har träffat en formell överenskommelse - att kommissionen är principiellt beredd att rätta sig efter dessa funderingar .
Beslut om detta kan dock inte fattas i och med denna förordning , utan det blir möjligt först inom ramen för den planerade revideringen av budgetplanen .
Genom förordningen , som sträcker sig över tiden 2000 till 2004 , får de båda förhandlande länderna rätt till tekniskt och finansiellt stöd för att införliva gemenskapens regelverk , för att kunna delta i gemenskapsprogram och särskilda inriktningar inom gemenskapen , liksom för att bygga ut kapaciteten inom sina förvaltningar och domstolar .
Av det planerade totalbeloppet på 95 miljoner euro tillfaller 57 miljoner euro Cypern och 38 miljoner euro Malta .
Vad gäller Cypern så omfattar förslaget till förordning även finansieringen av åtgärder som syftar till att stödja försoningen mellan de båda folkgrupperna , nämligen en tredjedel av det totala beloppet .
Jag skall från kommissionens sida se till att programplaneringen av anslagen görs i samklang med prioriteringarna inom partnerskapen för medlemskap redan under de kommande veckorna .
Och nu några korta kommentarer till hur Cypernfrågan har utvecklats efter Europeiska rådet i Helsingfors .
Jag kan helt och fullt sluta upp bakom vad statssekreterare Seixas de Costa har lagt fram på det portugisiska ordförandeskapets vägnar .
Vi har i denna fråga ett nära och bra samarbete .
Unionen har ju alltid sagt att medlemskapsförhandlingarna skall ha en positiv inverkan på lösningen av de politiska problemen på Cypern .
Vi har alltid varit införstådda med , och jag anser definitivt att det är riktigt , att förhandlingarna om lösningen på det politiska problemet skall föras under Förenta nationernas beskydd , och vi har alltid varit eniga om att lösningen fortsättningsvis skall vara en federation mellan två kommuner och två zoner som mål .
Det förblir Europeiska unionens mål att uppta ett förenat Cypern i unionen .
Rådet i Helsingfors har återigen betonat att en lösning på den politiska konflikten skulle underlätta medlemskap för Cypern i Europeiska unionen .
Emellertid , vilket ordförandeskapet redan har redogjort för , har rådet gett uttryck för att detta inte är några villkor för att förhandlingarna skall kunna avslutas .
Ifall en politisk lösning på Cypernfrågan inte har nåtts vid tidpunkten för de avslutade medlemskapsförhandlingarna skall rådet i betraktande av alla då relevanta faktorer fatta beslut om Cyperns inträde i unionen .
Så ser vårt politiska läge ut .
Europarådets beslut i Helsingfors om hur förbindelserna mellan Europeiska unionen och Turkiet skall gestaltas i framtiden har utvecklat stor dynamik .
Jag vill betona att det är ett flertal politiska processer som löper parallellt och är nära förbundna med varandra .
För det första gäller det förhållandet EU-Turkiet .
För det andra gäller det den fortsatta utvecklingen av de grekisk-turkiska förbindelserna , och det gäller fredsprocessen på Cypern .
Det har redan talats om ett window of opportunity , om möjligheternas fönster , som öppnar sig även till följd av den grekisk-turkiska avspänningen .
Vad kan vi då göra för att utnyttja detta möjligheternas fönster när det gäller problemet på Cypern ?
Jag tror att vi till en början måste välja en klok och återhållsam väg .
Om vi går för bryskt fram i den här frågan kommer vi att väcka förväntningar som inte kan infrias , utan jag är för ett förnuftigt agerande som får gå stegvis framåt och som är anpassat efter rådande situation .
Det första vi kan och vill göra är att förstärka dialogen och kommunikationen mellan de båda förbunden på Cypern .
Detta är en reflexion som understöds av våra grekiska och turkiska partner .
Vi vill alltså återuppliva de så kallade bikommunala aktiviteterna , och då framför allt bikommunala aktiviteter unga människor emellan .
Vi skall också i större utsträckning vinnlägga oss om att förbättra informationen om unionens mål till de turkcypriotiska förbunden .
Jag är fast övertygad om att en större förståelse av fördraget , ja större förståelse för vad Europeiska unionen egentligen är och vad den vill , att detta kan bidra till att undanröja rädsla och fördomar .
I mitten av mars kommer jag att resa till Cypern .
Mitt mål kommer att bli att bidra till att övertyga de båda förbunden om fördelen med ett nytt samarbete .
I den nya budgetförordningen har vi återigen avsatt medel för detta ändamål .
Det är inga oansenliga summor .
Det är mycket viktigt att vi vädjar till bägge sidor om att äntligen övervinna skuggorna från det förgångna och steg för steg utveckla en ny form för samarbete och slutligen för samlevnad .
Samtalen inom ramen för Förenta nationerna fördes i New York i december och i Genève i början av februari .
I maj kommer man att gå in i den kanske avgörande tredje rundan .
Förhandlingar skall i praktiken pågå ända tills en lösning har hittats , eller åtminstone tills man har gjort långtgående framsteg i de stora frågor som ordförandeskapet just har redogjort för .
Vad har då kommissionen för roll ?
Det är intressant att konstatera att alla inblandade i denna process anser att Europeiska unionens roll är central .
Alla inblandade i processen söker kontakt med och söker samarbete med oss .
Alla inblandade har klart för sig att fredsprocessen och tillämpningen av vårt gemensamma regelverk är oskiljaktigt förbundna med varandra och inte får råka i strid med varandra .
Jag måste säga att även jag sätter utomordentligt stort värde på samarbetet med Förenta nationernas generalsekreterare och dennes särskilda sändebud i ärendet och vågar påstå att det är ett samarbete som förlöper förtroendefullt och friktionsfritt .
Slutsatsen att det har blivit större dynamik i lösningen på Cypernfrågan efter Helsingfors är alltså berättigad .
Mycket längre än så vill jag för ögonblicket inte gå i min bedömning .
Unionens beslut att påbörja medlemskapsförhandlingarna och driva dem i jämn och rask takt , för att därmed även tjäna som katalysator i lösningen på det politiska problemet , är för mig fortfarande den rätta vägen .
Åtminstone ser jag inget på långa vägar förnuftigt alternativ till denna väg och kan därför bara säga att kommissionen kommer att hålla fast vid sin linje att ända till slutet av medlemsförhandlingarna även medverka till att det politiska problemet skall lösas samt att använda själva förhandlingarna om medlemskap som ett viktigt instrument i konfliktlösningen . .
( DE ) Herr talman , kära kolleger !
Jag tackar för de båda meddelandena och förklaringarna som kommissionär Verheugen just gav om förslaget till rådets förordning om genomförandet av åtgärder inom ramen för förberedelsestrategin .
Helt klart måste vi se Malta och Cypern som två kandidater som både politiskt sett och vad gäller förberedelsestrategin måste behandlas likvärdigt med de övriga 10 stater som det har inletts bilaterala förhandlingar med .
Säkerligen tvivlar ingen här i kammaren på att det skulle vara till utomordentligt stor hjälp om man lyckades finna en lösning på det cypriotiska problemet , och det råder heller ingen tvekan om att Europeiska unionen bör lämna sitt bidrag till detta .
Det vore en stor framgång om förhandlingarna kunde leda till att det blir ett enligt kommissionärens beskrivning förenat Cypern som går med i Europeiska unionen .
Å andra sidan måste vi naturligtvis också göra klart att det finns andra optioner , för att inte riskera att hamna i förlägenheter som i slutändan försätter oss i problem som driver hela utvidgningsfrågan till handlingsförlamning och blockad .
Redan de olika optionerna visar att detta kommer att bli ett av de kinkigaste problemen , om inte i slutändan det allra kinkigaste problemet i hela utvidgningen , där vi kanske kan vänta de största politiska svårigheterna .
Jag anser att det är utomordentligt viktigt att denna förberedelsestrategi nu förs på ett sådant sätt att dessa båda communities förenas redan på Cypern .
Cypern är , liksom Malta , på det hela taget ett relativt rikt land jämfört med övriga kandidatländer , men icke desto mindre måste det finnas ett visst mått av lika behandling .
På Cypern borde denna jämlika behandling också utnyttjas för att se till att den ekonomiska och sociala klyftan mellan den grekiska och den turkiska delen inte blir ännu större så att den ökade klyftan gör chanserna till ett enande ännu mindre .
Därför anser jag att denna förberedelsestrategi är alldeles särskilt betydelsefull .
Låt mig därför i all korthet ta upp de punkter som är viktiga i parlamentets ögon .
Jag vill tacka kommissionen för att man klart och tydligt har gått i ställning när det gäller klassificeringen i utgiftsområde B-7 , i den mån man så har kunnat i hittillsvarande beslutssituation .
Jag hoppas att även rådet kommer att ta samma steg och avge sin förklaring ; för Europaparlamentet står det nämligen utom allt tvivel att detta är en politisk fråga .
Det här ger överensstämmelse och rättvis placering i förberedelsestrategin , och samtidigt skall det garantera att siffrorna fram till år 2004 kan nämnas inalles så att budgetens tillförlitlighet , klarhet och sanningsenlighet tryggas även i det här fallet .
Som det har skötts hittills får man inte ihop det med ett normalt budgetförfarande .
Jag anser att det är viktigt att säga att Europaparlamentet ändå har medverkat positivt för i år eftersom vi inte vill att dessa länder skall få några nackdelar , varför vi var beredda att fatta de nödvändiga besluten för budget 2000 , men det kan också bara gälla just för i år .
Därför är det av vikt att ordförandeskapet i samband med överläggningarna kring betänkandet författar motsvarande meddelande som gör det möjligt för oss att ta upp frågan i en ordnad process på det att detta i mina ögon så onödiga gräl kan få ett slut .
Jag har stor förståelse för att det kan uppstå matematiska problem här på grund av Agenda 2000 och det kapital som må stå till förfogande .
Jag vill också klart och tydligt säga att man kanske rentav kan förhandla om siffran 130 miljoner , som nämns i mitt betänkande .
Det har lämnats in ett ändringsförslag från kammaren till i morgon , vilket utgår från ett annat belopp , i synnerhet som dessa länder , som jag sade , ju har en relativt hög utvecklingsnivå .
Likväl måste det finnas en säkerhet i dessa länder för den närmaste förutsebara tiden , de måste veta vad de faktiskt har att vänta sig , och detta måste också avspegla sig i planeringen i Europaparlamentet som en del av budgetmyndigheten .
Herr rådsordförande , jag vet att ni alltid har den goda viljan när det gäller samarbetet med Europaparlamentet .
Jag hoppas att så är fallet med rådet som helhet samt att ni skall kunna ge oss de rätta svaren på dessa frågor . - ( EL ) Herr talman !
Vi har hört rådets och kommissionens uttalanden , och jag skulle vilja göra följande kommentarer : Herr rådsordförande !
Jag förstår den försiktighet med vilken ni bemöter ämnet och era ansträngningar i kontakterna med den turkcypriotiska sidan , men kanske skulle det vara tydligare och korrektare om den vokabulär som ni använder inte gav upphov till misstankar om att ni kanske eftersträvar något slags indirekt erkännande , trots att ni har betonat att så inte är fallet .
Till exempel skulle jag inte säga Nicosias regering .
Det rör sig om den cypriotiska regeringen , herr rådsordförande , det rör sig inte om Nicosias regering .
Denna regering har föreslagit ett tillvägagångssätt som gör att den turkcypriotiska sidan kan delta , och jag anser att det rätta för rådet och kommissionen att göra är att trycka på den turkcypriotiska sidan att delta institutionellt inom ramen för de förhandlingar som förs av Republiken Cypern .
Å andra sidan väcker det sätt som frågan om slutande av protokollen och föranslutningsstrategin hittills har behandlats på vissa tvivel .
Jag förstår inte varför det bör göras ett undantag för de två små länderna , eller varför det behövdes en konflikt mellan institutionerna eller påtryckningar från parlamentet för att få in medlen i kapitel 7 om föranslutningsstrategin .
Bör verkligen Europeiska unionen behandla två små länder i utkanten av unionen på detta sätt ?
Det rör sig ju om länder som unionen behöver , men som även har allt det som behövs för att kunna fungera i unionen och som anses redan skulle kunna delta i den ekonomiska och monetära unionen ?
Som kommissionären sade - och jag instämmer med honom - är det fråga om ett politiskt beslut .
Och det rör sig om ett litet politiskt beslut , herr rådsordförande , med tanke på de stora fördelarna , och framför allt med tanke på den hjälp det skulle kunna ge de två folkgrupperna att verkligen utgöra en stat , och förbindelserna måste återupptas - ­ för det har tidigare funnits förbindelser mellan de två grupperna - - , och Republiken Cypern måste verkligen befrias från ockupationsstyrkorna .
Herr talman , kära kolleger !
Inom ramen för samrådsförfarandet har vi behandlat ett förslag till rådets förordning , om genomförande av åtgärder inom ramen för en strategi inför anslutningen för Cypern och Malta .
Detta förslag påminner om dem som har lagts fram för de övriga kandidatländerna , och när det väl genomförs kommer det att ersätta de finansprotokoll som nu har upphört att gälla .
Instrumenten inför anslutningen syftar till att ge ett tekniskt och finansiellt bidrag till kandidatländernas ansträngningar för att uppfylla kraven i gemenskapens regelverk .
Kommissionens analys har faktiskt visat att Cypern och Malta - trots att de ingår i Världsbankens kategori med höginkomstländer - uppvisar samma svårigheter som länderna i Central- och Östeuropa att införliva gemenskapsrätten , på grund av att de saknar en tillräcklig administrativ och juridisk kapacitet .
När det utmärkta betänkandet av Brok behandlades i utskottet , klargjordes det att dessa två länder också kan komma ifråga för stöd enligt budgetposten Meda , för övergripande åtgärder av regionalt intresse .
Jag skulle vilja be kommissionären att bekräfta detta tydligt .
När det gäller Cypern måste man precisera att en del av det tekniska och finansiella stöd som instrumenten föreskriver är avsett för ett närmande mellan den grekiska och den turkiska gemenskapen och en definitiv lösning på problemet med öns delning .
Rådets och kommissionens uttalanden om den cypriotiska frågan var därför särskilt lämpliga , och jag vill tacka rådets ordförande och kommissionär Verheugen .
Sedan den 4 juli 1990 , då Cypern lämnade in sin ansökan om medlemskap , har Europaparlamentet antagit en mängd resolutioner för att kräva en politisk lösning i enlighet med internationell rätt och de tillämpliga resolutionerna från Förenta nationernas säkerhetsråd .
I april 1999 upprepade parlamentet sin ståndpunkt , dvs. att Cyperns anslutning till EU skall komma hela ön till del samt underlätta en politisk lösning , men att det sistnämnda inte skall utgöra ett villkor för ett medlemskap .
Med andra ord skall en politisk lösning inte hålla EU-anslutningen som gisslan .
De två processerna är två separata processer .
Denna otvetydiga ståndpunkt från kammarens sida har väckt en del kontroverser .
Vi skall alltså glädja oss åt att Europeiska rådet i Helsingfors satte stopp för spekulationerna genom att slå fast följande i slutsatserna : " har man inte nått fram till en lösning när medlemskapsförhandlingarna är avslutade , kommer rådet att fatta beslut om ett medlemskap utan att det ovannämnda utgör en nödvändig förutsättning " .
Eftersom situationen är klar , får vi nu hoppas på att förbättrade förbindelser mellan Europeiska unionen och Turkiet och bättre grekisk-turkiska förbindelser får en gynnsam inverkan på det turkcypriotiska samhället , och att turkcyprioterna inte längre kommer att vägra att skicka företrädare till medlemskapsförhandlingarna .
Det faktum att dessa företrädare närvarar skulle på intet sätt avgöra den definitiva politiska lösningen .
Snarare tvärtom .
Detta gör att samtliga parters intressen kan värderas , vid ett ögonblick då Cypern infogas i Europeiska unionen och därmed gör sig berett att ta ett avgörande steg i sin historia .
Herr talman !
Jag vill också ansluta mig till föredragandenas glädje över att man nu ser bättre möjligheter för att komma vidare när det gäller utvecklingen på Cypern , i takt med att förhållandet mellan Turkiet och EU och mellan Turkiet och Grekland har blivit bättre .
Men jag tycker också att EU skall ge ett konstruktivt bidrag .
Jag tycker också - vilket redan nämnts - att det finns vissa problem med budgetförordningen som vi måste lösa .
Det handlar ju om ett föranslutningsstöd och det hör hemma i utgiftsområde sju .
I fjol accepterade parlamentet undantagsvis att pengarna till dessa utgifter placerades i utgiftsområde fyra och därmed behandlas de två ansökarländerna inte likvärdigt med ansökarländerna från Central- och Östeuropa , och så skall ju ske enligt förklaringarna från toppmötet i Helsingfors .
Det skall alltså avsättas medel i utgiftsområde sju , där det skall ske en revidering av budgetplanerna .
Detta är den springande punkten .
Huvudsaken är att pengarna till Cyperns och Maltas föranslutningsstöd hämtas från utgiftsområde sju och att det sker en revidering av budgetplanerna , därför om rådet inte accepterar detta agerar det ju i realiteten i strid mot sina egna beslut i Helsingfors i december .
Vad gäller det belopp som anges i Brokbetänkandet , 130 miljoner euro , vill jag också på den liberala gruppens vägnar säga att vi måste komma fram till ett belopp , vi måste förhandla oss fram till beloppets storlek .
Det viktigaste är att ett flerårigt program säkerställs och i den rätta utgiftsområdet , så att Cypern och Malta kan börja planera .
Herr talman !
Gruppen De Gröna / Europeiska fria alliansen stöder det beslut som rådet fattade i Helsingfors , enligt vilket en lösning på konflikten inte får utgöra en förutsättning för Cyperns medlemskap .
Regeringen på Cypern måste utsättas för ett hårt tryck , men viljan hos en majoritet av befolkningen får inte utsättas för blackmail , utpressning , från en del av befolkningen , eftersom vi anser att man kan hysa starka tvivel när det gäller regeringens representativitet på den delen av ön .
Det är uppenbart att detta möjligheternas fönster - " la janela de oportunidades " , som ordförandeskapet uttryckte saken - måste utnyttjas maximalt .
Jag är även övertygad om , trots att de turkisk-grekiska förbindelserna har förbättrats , att detta inte räcker .
Lösningen på Cypernkonflikten står framför allt att finna i en förbättring av förbindelserna mellan de båda samhällena , i väntan på - och vi hoppas att väntan inte blir för lång - en federation .
Vi måste framför allt verka för att man löser frågan om fri rörlighet , problemet med demilitariseringen och att vapnen försvinner från ön .
Europeiska unionen borde spela en mer framträdande roll , utöver det ekonomiska stödet - som i och för sig är viktigt - som garant för och främjare av kontakter mellan de olika samhällena och inrätta fora och program för confidence building .
Låt mig säga att i detta ögonblick känner jag starkt saknaden efter Alex Langer i parlamentet , Alex Langer som var en fredsbyggare och ett föredöme för oss alla när det gäller hur man bygger upp en samexistens mellan olika folk .
Herr talman !
Försöken att frammana en dialog mellan de två cypriotiska parterna under FN : s beskydd erinrar oss om att ockupationen fortfarande pågår 26 år efter den turkiska arméns invasion av ön ; på 40 procent av territoriet finns 35 000 soldater , tung militär utrustning och 50 000 kolonisatörer , vilket strider fullständigt med resolutionerna från Förenta nationernas säkerhetsråd i den här frågan .
Vad kan Europeiska unionen göra i det här sammanhanget , något som inte utgör en inblandning i frågor som endast cyprioterna kan avgöra , men som kan främja strävan efter en rättvis och bestående lösning på detta dramatiska problem , ett problem som drabbar ett land som i nästan 30 år har haft förbindelser med Europeiska gemenskapen och som är kallat att integreras i unionen under de kommande åren ?
Jag har hört uttalanden och uppfattat en något tvetydig tystnad , bland annat från rådets sida , och det är något som i mina ögon borde klargöras .
Det första som åligger oss tror jag är att erinra om den viktigaste referensen i den här frågan för hela världssamfundet - Förenta nationernas resolutioner .
Enligt säkerhetsrådet bör en lösning på det cypriotiska problemet bestå i en federation med två områden , två samhällen , med andra ord - Verheugen anspelade på detta - en enhetsstat som inbegriper två lokala administrationer som skall företräda de två samhällena .
Suveräniteten , statusen av internationell person och medborgarskapet skall vara enhetligt och denna stat bör demilitariseras .
På så sätt markerar världssamfundet att det inte accepterar ett fullbordat faktum uppnått med våld .
För det andra tror jag att Europeiska unionen vinner på att så långt det är möjligt begränsa tolkningsmöjligheterna av den ståndpunkt som fastställdes av Europeiska rådet i Helsingfors .
Lösningen på det cypriotiska problemet får inte vara en nödvändig förutsättning för Cyperns anslutning till unionen , vilket Poos erinrade om .
Det motsatta alternativet skulle innebära att Turkiet anförtros en sorts vetorätt i fråga om Cyperns anslutning till Europeiska unionen , vilket självklart inte är godtagbart .
För det tredje slutligen : Europeiska rådets ståndpunkt från Helsingfors får i gengäld inte leda till att vi dämpar våra ansträngningar för att lösa det cypriotiska problemet innan landet skall träda in i unionen .
Ur den synvinkeln skänker det andra beslutet från Helsingfors ett nytt ansvar , och samtidigt nya möjligheter , till de 15 EU-medlemmarna - dvs. erkännandet av Turkiets ansökan om medlemskap i unionen .
EU : s dialog med Ankara kan och bör , i mina ögon , avse den fast beslutna viljan att få Turkiet att visa en konstruktiv attityd gentemot dialogen mellan de två cypriotiska samhällena och därmed en respekt för internationell legalitet , vilket skulle kunna mynna ut i ett återförenat Cypern och fred i östra Medelhavsregionen .
Herr talman !
I fråga om vikten av ekonomisk hjälp till Cypern och Malta förekommer inga större meningsskiljaktigheter .
Den stora frågan är snarare under vilket budgetområde denna hjälp skall finansieras .
Rådet och kommissionen föreslår att låta protokollen falla under utgiftsområde 4 .
Det överensstämmer med parlamentets budgetbeslut i december .
Föredraganden återkommer till detta och föreslår nu att föra in Cypern och Malta utgiftsområde 7 .
Budgetutskottet föreslår till och med att godkännandet av Brokbetänkandet skall skjutas upp tills rådet kommer med ett löfte om att höja finansieringsramen för utgiftsområde 7 .
Det är en ytterst riskabel strategi .
Utan omröstning i parlamentet kan ju inte finansprotokollen starta .
På det sättet går det politiska spelet mellan rådet och parlamentet om storleken för ramarna ut över Cypern och Malta .
Dessutom , vad är finansieringsramar värda om de höjs vid varje ny åtgärd ?
Jag skulle därför vilja förespråka att låta de 15 miljonerna euro i enlighet med kommissionens förslag falla under utgiftsområde 4 .
När det gäller krediterna för de kommande åren kan en flerårsbudget från kommissionen , senare under året , ge närmare besked .
Herr talman !
Runt om i världen arbetar man för att lösa långvariga konflikter och föra samman folkgrupper som har delats av historien och av gammalt fiendskap och hat mellan grupperna .
Det är nu vi måste ägna vår tid och kraft åt att hjälpa cyprioter från båda sidor av den " gröna linjen " att finna en lösning på en konflikt som har varat allt för länge .
Vi vet alla att det krävs särskild omsorg för att säkerställa att Cypern framgångsrikt förs in i Europeiska unionen , och de beslut som fattades i Helsingfors ger ytterligare en dimension till denna debatt , med godkännandet av Turkiet som ett kandidatland .
Jag hoppas att de beslut som fattades i Helsingfors leder till framsteg i Cypernfrågan .
Jag hoppas att detta signalerar en ny era av hopp för Cypern .
Jag hoppas att Turkiet börjar spela en konstruktiv roll Cypernfrågan .
Jag blir mycket glad av att höra de stödjande orden från rådet och kommissionen för FN och för organisationens arbete med att uppmuntra närhetsamtal mellan de två folkgrupperna i syfte att uppmuntra försoning och återuppbyggnad av förtroende mellan de två folkgrupperna på Cypern .
Jag välkomnar kommissionens stöd för detta två zoners och två gruppers federala Cypern som FN har arbetat för så länge och som både den grekcypriotiska sidan och den turkcypriotiska sidan borde arbeta hårt för att förverkliga .
Jag välkomnar den förnyade värmen i förbindelserna mellan den grekiska regeringen och den turkiska regeringen .
Jag hoppas att den har en uppmuntrande effekt på Cypernsamtalen .
Jag hoppas att de anslutningsmedel som finns tillgängliga för att hjälpa Cypern delvis används till att främja försoningen och förtroendeuppbyggnaden samt att båda sidor av de delade folkgrupperna på Cypern godtar och använder dessa medel i samma anda som de ges .
Vi bör alla , i alla de europeiska institutionerna - i parlamentet , rådet och kommissionen - , göra vårt bästa för att hjälpa Cypern i dess strävan att nå en fredlig lösning som för samman dessa två folkgrupper , vilka har varit delade under allt för många år .
Herr talman , kära kolleger !
Först vill jag tacka ordförandeskapet , tjänstgörande rådsordförande Seixas da Costa och kommissionär Verheugen för redogörelserna om Cypern .
Det gläder mig mycket att bägge två har understrukit att Europeiska unionen tänker arbeta hårdare för att få en lösning på Cypernfrågan .
För vi alla vet att det är oacceptabelt att ön har varit delad sedan 1974 , att runt 38 procent av Cypern har varit ockuperat av Turkiet i mer än 26 år .
I det förgångna har alla försök att finna en fredlig lösning på Cyperns problem strandat på den turkiska sidans orubbliga hållning samt på den turkcypriotiska ledningen .
Men jag tror , vilket också blev tydligt i era ord , att vi nu i början av detta år 2000 möjligtvis har fått en ny situation och att vi eventuellt har nya chanser .
För det första ser vi Förenta nationernas nya åtgärder , vilket redan har diskuterats ; vi ser nya åtgärder från USA : s regering , vi ser ett tydligt närmande mellan Turkiet och Grekland .
Men i synnerhet efter rådets beslut i Helsingfors tror jag att man kan vänta sig ett genombrott .
I Helsingfors upptog unionen Turkiet i kretsen av kandidatländer .
Samtidigt beslutades det att lösningen på Cypernfrågan inte är något villkor för att Cypern skall kunna gå med i unionen , vilket egentligen - kollegan Poos poängterar detta - var ett klart ställningstagande från unionen och från parlamentet , vilket också har bekräftats i olika resolutioner .
Turkiet vet alltså utan tvivel från Helsingfors att de inte har någon vetorätt i fråga om Cyperns medlemskap och att deras fortsatta fördjupande av förbindelserna till Europeiska unionen är nära förbundet med lösningen på Cypernfrågan .
Därför får man verkligen hoppas att några kloka politiker i Ankara ser den chans som ett slut på den turkiska ockupationen av Cypern innebär för Turkiet självt .
Jag hoppas verkligen att - som det har sagts här - detta chansernas eller möjligheternas fönster verkligen ställs på vid gavel och att även företrädare för rådet och kommissionen arbetar vidare i denna riktning i Ankara .
Men i motsats till Frassoni anser jag inte att Cypernfrågan endast är en fråga för folkgemenskaperna , utan i allt väsentligt en fråga för den turkiska politiken .
Jag tror att vi kan utgå ifrån att Cyperns process mot ett medlemskap i EU inte kan avbrytas .
Och vi hoppas alla att det skall bli ett förenat Cypern som går med .
Därför har jag en fråga om ett klarläggande till er , herr ordförande : Ni talade om deltagandet från den turkcypriotiska sidan .
Finns det någon form av signaler om att den turkcypriotiska sidan kommer att gå med på den cypriotiska regeringens eller Europeiska kommissionens anbud och att man kommer att vilja anta erbjudandet om att delta i samtalen ?
Vad gäller den andra punkten : Det gläder mig mycket att vi utifrån Brokbetänkandet - och hjärtligt tack för betänkandet , herr föredragande - denna vecka också tar itu med de finansiella aspekterna på förberedelsestrategin för Cypern och Malta .
För det krävs absolut att det ges finansiell hjälp för anpassningen till det gemensamma regelverket när finansprotokollet för Cypern och Malta har löpt ut .
De två länderna hör helt säkert inte till de fattigaste kandidatländerna .
Men anpassningsåtgärderna är omfattande även för Cypern och Malta .
För anpassningsåtgärderna mellan 1999 och 2002 räknar Cypern med utgifter på runt 850 miljoner euro , vilket motsvarar knappt 12 procent av den egna bruttonationalprodukten .
Därför har utskottet för utrikesfrågor talat för en ökning av det planerade beloppet på 95 miljoner euro .
Och jag hoppas verkligen att vi faktiskt skall ha möjlighet att öka på beloppet .
För cyprioternas skull , de grekiska liksom de turkiska , får man hoppas att väsentligt kapital kan flyta in till de planerade åtgärderna för ett bikommunalt samarbete , vilket kommissionär Verheugen ju nämnde , i syfte att få de båda folkgrupperna att närma sig varandra igen .
Jag har en sista fråga till kommissionär Verheugen : Har ni fått några signaler på att bikommunala kontakter på Cypern har bättre förutsättningar nu än efter Luxemburg ?
Där försvann ju möjligheterna i och med förbudet från Denktash .
Herr talman , kära kolleger , bäste herr rådsordförande , bäste kommissionär Verheugen !
Förordningen för medlemskapsstöden är inte direkt ett lysande exempel på samstämmigheten i kommissionens arbete .
Detta hopkok av hjälpkonstruktioner ger snarare ett intryck av dilettanteri .
Det gäller såväl den innehållsliga utformningen som den finanstekniska aspekten .
Därmed , anser jag , kan vi svårligen presentera unionens medlemskapsåtgärder för medborgarna på Cypern och Malta som ett bevis på att det lönar sig att gå med .
Vaclav Havel har i dag med rätta sagt att Europeiska unionens politiska kvalitet bedöms efter vad den enskilda människan får ut .
Ur det medborgerliga samhällets synvinkel är det vad en förordning ger som är det avgörande .
Med den här förordningen uppnår man inte precis det perfekta .
Den innehåller artiklar som inte baseras på självbestämmande och den är provisorisk , och det är ingenting att briljera med .
Kvalitén på bidragshjälp mäts enligt följande måttstock : Är den decentralistisk , är den genomblickbar , står den nära medborgarna samt fungerar den ?
Icke desto mindre , för den delade ön Cypern är denna föranslutningsstrategi på det hela taget förenad med en stor politisk utmaning .
Som jag ser det består Europeiska unionens uppgift i att utnyttja alla verktyg , även detta , för att bidra till en politisk konfliktlösning på ön .
Här måste jag säga att just Europaparlamentets ändringsförslag är mycket viktigt för mig .
Även från kommissionens och rådets sida hålls det i dag mycket hoppingivande tal .
Jag är mycket , mycket glad att vi har en och samma inriktning här .
För mig är preferensoptionen verkligen att Cypern i och med en fredslösning i landet tas upp i Europeiska unionen .
Herr rådsordförande , herr kommissionär !
I Greklands kommunistpartis ögon är Cyperns huvudsakliga problem inte dess anslutning till Europeiska unionen utan den turkiska ockupationen av 40 procent av Cyperns yta , som har pågått i 26 år .
Det cypriotiska folkets framtid går genom detta lilla lands enande , oberoende av varje cypriots nationella ursprung .
Den enda godtagbara lösningen som garanterar framtiden och som inte kommer att erbjuda några möjligheter till utländsk inblandning , som den typ av inblandning som har framkallat den senaste femtioårsperiodens alla problem , är ett enat och federalt Cypern , i enlighet med resolutionerna från FN : s säkerhetsråd .
Nyckeln till lösningen på Cypernfrågan finns i händerna på den turkiska regeringen , som stöder och uppmuntrar den turkcypriotiske ledarens , Rauf Denktash , kompromisslöshet .
Europeiska unionen , med sitt spelade intresse för frihet och mänskliga rättigheter , har å sin sida aldrig låtit sig beröras av det cypriotiska folkets tragedi , av problemet med de grekcypriotiska och turkcypriotiska flyktingarna , av den våldsamma förändringen i befolkningssammansättningen på norra Cypern , av Turkiets kraftiga utplacering av bosättare på de ockuperade områdena .
Till och med här i denna sal talade rådets ordförande om Cyperns norra del och inte om de ockuperade områdena .
Beslutet i Helsingfors nyligen att ge Turkiet status som kandidatland , utan att landet har gjort den minsta eftergift i frågan om Cyperns ockupation , som till exempel att minska sin militära närvaro på ön eller att återlämna Ammokosto , uppmuntrar utan tvekan den turkiska kompromisslösheten .
Uttalandena av den turkiske premiärministern , Bülent Ecevit , omedelbart efter Helsingforsmötet om att Cypernproblemet löstes 1974 är ingen tillfällighet .
Att uppmuntra den turkiska kompromisslösheten gör det naturligtvis inte lättare att föra de två folkgrupperna närmare varandra i de nära förestående samtalen som kommer att föras under FN : s generalsekreterares beskydd .
På sin väg mot anslutning har Cyperns folk redan förlorat mycket , men det kommer att förlora ännu mer .
Genomförandet av gemenskapens regelverk har skapat allvarliga problem i den cypriotiska ekonomin , särskilt inom jordbruket , det innebär krav på att den offentliga sektorn skall säljas ut och det medför att det utvecklade sociala solidaritetssystem som finns i landet rivs ned och förstörs .
Herr talman !
Ursäkta mig , men det gjordes ett litet översättningsmisstag i den franska hytten , vilket gäller Alyssandrakis ord , det känsligaste ordet i hela debatten .
Jag vill inte att det skall råda tvivel på denna punkt .
Den franska översättningen fick Alyssandrakis att säga att " en konfederal lösning är den bästa " .
Det är uppenbart att Alyssandrakis sade : " en f e d e r a l lösning är den bästa " .
Det är mycket , mycket viktigt att detta klargörs , herr talman .
Stort tack för klarläggandet , herr Wurtz .
Herr talman !
Malta och Cypern skiljer sig mycket från länderna på Europas fastland .
Särskilt malteserna har varit mycket duktiga på att överleva under fientliga geografiska och geopolitiska förhållanden .
Deras framgång har till stor del vilat på deras företagsamhet , deras dynamiska kraft och deras flexibilitet .
Malta har en sjudande lätt och tung industri , en växande marknad för finansiella tjänster , ett bra jordbruk , utmärkt turism och ett häpnadsväckande urval arbetstillfällen - och allt detta på en ö som så gott som helt saknar naturresurser .
Jag är därför övertygad om att en ö som Malta , med sin befolkning på 340 000 , inte kan anpassa sig till rigiditeten i de ekonomiska och rättsliga strukturerna från fastlandet , som har en befolkning som är tusen gånger större .
När jag betraktar det föreslagna instrumentet , ser jag följaktligen inte en åtgärd som skall föra två folk in i moder Europas hägn .
Situationen är mer att likna vid ett svart hål i rymden , som suger till sig massa med en sådan kraft att inte ens ljuset undkommer .
Vi borde inte muta dessa ömänniskor till att samarbeta till sin egen undergång , genom att ge dem pengar för att ta till sig lagar som är lika främmande för deras kultur som ett svart hål är för moder jord .
EU borde lämna Cypern och Malta i fred .
I mina ögon verkar det som att de enda människorna på Malta som vill detta är den politiska klassen , och jag skall hålla tummarna för att det maltesiska folket återigen kommer att stå som vinnare .
Herr talman !
Att döma av inläggen från kollegerna i detta parlament , från alla sidor , är detta en av de få gånger som det råder en mycket stor enighet om Cypernfrågan , liksom naturligtvis om anslutningsförfarandet för Cypern och Malta .
Det betyder att det finns ett gemensamt medvetande hos oss alla om Cyperns , som det heter , politiska problem .
Samtidigt innebär det emellertid att ett mycket stort tryck sätts på både rådet och kommissionen att låta denna samstämmighet , som är ett uttryck för Europas partiers och alla folks vilja , utgöra utgångspunkt för deras eget sätt att angripa problemet .
Mina damer och herrar !
Helsingforsmötet var ett historiskt möte , en historisk vändpunkt , en ny historisk referenspunkt .
Om några personer av någon som helst anledning skulle anse att den balans som nåddes där utgör en utgångspunkt för nya förhandlingar någon annanstans , om några personer med sin egen hållning skulle destabilisera denna helhet av fakta och balans , skulle de begå ett tragiskt misstag .
Omständigheterna är mogna .
Vad som krävs av Europeiska unionen , av rådet , av alla , är en lugn beslutsamhet , en lugn beslutsamhet att utan knep och manövrer fortsätta anslutningsförhandlingarna med både Cypern och Malta - som när allt kommer omkring är de mest mogna av alla ansökarländerna - , så att denna beslutsamhet kan fungera som en referenspunkt för varje sida som kan ha en annan åsikt än den som vi alla instämmer i .
Broks betänkande är ett bra verktyg i denna riktning , och det faktum att betänkandet på grund av att diskussionen är gemensam täcks in politiskt av rådets och kommissionens politiska anföranden är faktiskt litet beklagligt , och vi kan följaktligen inte säga fler saker om detta goda betänkande .
Under alla omständigheter befinner sig utvecklingen i era egna händer .
Utvecklingen befinner sig i våra egna händer , i så måtto att vi utrustar er med beslut , i så måtto att vi utrustar er med möjligheter .
Angående Broks betänkande , är Cypern och Malta de sista öarna i Medelhavet , och , om jag inte bedrar mig , i hela Europa , som ännu inte har anslutits till Europeiska unionen .
Detta har ett symboliskt värde , eftersom Medelhavet och dess öar - jag kommer själv från en ö - är den region som de människor som kommer från norra Europa för att fira sin sommarsemester och de människor som bor där huvudsakligen kommer i kontakt med .
Ur den synvinkeln är Afrodites ö , som Cypern kallas , och piraternas , som vi öbor med stor kärlek kallar maltesarna , ö två diamanter som snabbt måste införlivas i Europeiska unionen .
De har väl fungerande ekonomier , de har goda ekonomiska förbindelser , och de utgör , när allt kommer omkring , ett område där Europeiska unionens politiska vilja skall sättas på prov .
Avslutningsvis vill jag , då jag inte tycker att jag behöver bli långrandig , eftersom jag har noterat den enighet som råder i denna fråga , bara komma med en liten kommentar till rådsordföranden : Jag tycker att det på något ställe i hans anförande fanns vissa besynnerligheter , jag hoppas att det var översättningen som var felaktig , och jag hoppas att han tar upp saken i sin sammanfattning .
Herr talman !
Jag är den siste talaren , och därför skulle jag vilja ställa en fråga till Seixas da Costa och Verheugen , om Verheugen sätter på sig hörlurarna och om han är intresserad av att lyssna till alla talare .
Det handlar om två folkgrupper , men det handlar inte i första hand om två folkgrupper .
Som många talare har påpekat , rör det sig här om en ockupation .
Ett av Europeiska unionens kandidatländer - Turkiet - ockuperar en del av ett annat av Europeiska unionens kandidatländers yta .
Det finns där en militär styrka på 40 000 man , och Berlinmuren finns i dag i Leukosia .
Vi kan inte säga vad som kommer att hända - förutom i samtalen mellan Denktash och Republiken Cyperns president .
Den fråga som jag vill ställa framför allt till Seixas da Costa , men även till Verheugen , är följande : Vilka frågor tar rådet upp med den turkiska regeringen , med anledning av associeringsrådet , angående detta ?
Vilka frågor kommer rådet att ta upp angående trupptillbakadraganden , men även angående den turkiska regeringens bidrag till en lösning på Cypernfrågan ?
Jag vill påminna om att den turkiska regeringen , efter ett beslut nyligen i Europadomstolen för de mänskliga rättigheterna i Strasbourg , fälldes för expropriering av grekisk egendom .
Inte Denktash .
Inte något juridiskt diffust som " Turkiska republiken på norra Cypern " , utan den turkiska regeringen .
Jag frågar er : vilka frågor kommer med anledning av associeringsrådet att tas upp angående Turkiets bidrag till att finna en lösning på Cypernfrågan ? .
( PT ) Herr talman , ärade kollegor !
Jag har uppmärksamt lyssnat på vad som sagts , särskilt det som så emotionellt sades om Cypern , nämligen att för att försvara det som i dag är lag i Cypern så måste Europeiska unionen erkänna just de resolutioner som faller under Förenta nationernas säkerhetsråd i den här frågan .
Om detta finns ingen som helst tvetydig tystnad från rådets sida .
Rådet tar på sig allt ansvar vad gäller tolkningen av situationen i Cypern .
Det var för övrigt den situationen och den tolkningen som fick rådet att anta det beslut som antogs i Luxemburg i slutet av 1997 när man beslöt att ta de första stegen för en anslutning av Republiken Cypern till Europeiska unionen .
Jag vill så gärna försöka få ledamöterna att förstå att oberoende av de mer eller mindre emotionella ståndpunkterna i den här frågan så kräver de dagliga internationella förhandlingarna normalt sett att regeringarna , och när jag säger regeringar så menar jag alla , intar en mera flexibel inställning .
Vi behöver faktiskt ståndpunkter av en mera emotionell natur för att se till att vi förstår att alla de här frågorna rör människor , men vi måste också veta att det är genom förnuftiga politiska ståndpunkter och förhandlingsflexibilitet som man lyckas nå lösningar som kan se bortom de stora meningsskiljaktigheterna , vilka i grund och botten är orsak till många historiska tragedier .
Oavsett vem som är skyldig - och vi är inte här för att föra register över de skyldiga , Förenta nationernas resolutioner i den här frågan är tydliga - så menar jag att vi utan sinnesrörelse och på ett mera rationellt sätt bör ta tillvara de möjligheter som den nya situationen ger vid handen .
Europeiska rådet i Helsingfors hade mod att fatta vissa beslut , och jag tror att en del av de här besluten redan har börjat öppna de dörrar som går att öppna , som jag inledningsvis sade om möjligheternas dörr .
Konkreta resultat kan vi inte nå genom att utnyttja konflikter , inte i det här skedet av förhandlingarna , eftersom det är ett mycket känsligt skede .
Det är genom diskret arbete , genom att stödja sändebudet för Förenta nationernas generalsekreterare i hans uppdrag , det är så som vi måste fortsätta att arbeta .
Ärade kollegor , Europeiska unionen har intagit fel ståndpunkt i den här frågan , och det är förmodligen meningslöst att gå igenom de uttalanden som eventuellt kan finnas i rådets tal eller i vilken annan åsiktsförklaring som helst .
Vi är inte ute efter det politiskt korrekta i det här parlamentet .
Vi är ute efter det som internationellt sett är rättvist , vi är ute efter gemensamma ståndpunkter , ståndpunkter som allt efter som har definierats av rådet , som är hållbara och som Europeiska kommissionen omsorgsfullt , uppmärksamt och på ett pragmatiskt sätt också har följt .
När man säger att norra Cypern inför en eventuell framtida anslutning av Republiken Cypern till Europeiska unionen måste få ta del av informationsutbytet , så måste vi vara medvetna om att det vi håller på med är att försöka finna praktiska alternativ för att klara av de hinder som ligger i vägen för en politisk resolution .
Vi försöker inte hitta på några undanflykter och vi försöker inte , genom praktiska lösningar eller på annat sätt , finna något som kan vara ett erkännande av politisk natur .
Enligt min mening gav rådet i Europeiska unionen allteftersom klara besked om att detta inte är deras ståndpunkt .
Rådet har antagit besluten med stor ansvarskänsla .
Det som hände i Helsingfors är som vi ser det självklart .
Det sätt som vi har varit i förbindelse med Republiken Cypern under anslutningsförfarandet är något som till och med de inhemska myndigheterna i Republiken Cypern ser som mycket positivt .
Det är ingen mening att göra eller försöka göra en andra tolkning av våra avsikter .
Herr talman , mina damer och herrar !
Jag vill tacka så hjärtligt för debatten som jag på det stora hela uppfattar som en uppmuntrande och stödjande debatt som visar att det i kammaren råder stor enighet i medlemsstaternas politik och även i kommissionens .
Men jag vill gärna komma med ytterligare ett par klarlägganden som har efterfrågats .
För det första det som gäller ärendet med rubrikerna 4 och 7 .
Det är mycket enkelt : I Berlin har det , i samband med det stora Agenda 2000-paketet , upprättats en särskild rubrik för de öst- och centraleuropeiska kandidatländer som befinner sig i en omvandlingsprocess , nämligen just den berömda rubrik 7 , och då endast för dessa länder .
Malta , Cypern och Turkiet räknade man inte med då .
Fru Schroedter betecknade detta som en brist på samstämmighet .
Kanske skulle ni någon gång behöva fråga den dåvarande rådsordföranden , som ju inte är er så främmande , om hur denna som ni förmodar brist på samstämmighet har uppstått .
Även jag var i någon mån inblandad .
Jag tror inte att det är så , utan orsaken till beslutet var att man ville ha ett särskilt instrument för de öst- och centraleuropeiska staterna , vilka det ställs andra krav på under medlemskapsprocessen än på Malta och Cypern .
Likväl har jag sagt att jag förstår de argument som framförs här , och kommissionen kommer att bemöda sig om att ta hänsyn till dessa önskemål , men när det nu är Agenda 2000 och den budgetplanen det handlar om kan vi inte göra så utan att ändra i denna budgetplan .
Hittills har detta förstås inte alls varit möjligt .
Ett klarläggande : Om vi flyttar över det från rubrik 4 till rubrik 7 påverkas inte helhetsbalansen i budgeten .
Om vi gör det skulle rubrik 7 ökas och rubrik 4 minskas med motsvarande belopp .
Föreställningen om att man däremot skulle kunna lägga till det under rubrik 7 och låta rubrik 4 stå som den är går inte att genomföra .
Inte heller parlamentet kan göra av med pengar som man inte har , åtminstone inte så länge vi saknar en press stående i källaren att trycka eurosedlar med !
När det då gäller fredsprocessen på Cypern och kopplingen till medlemskapsförhandlingarna så vill jag upprepa att det alltid har varit så att medlemskapsförhandlingarna har stått i direkt samband med processen .
Det har alltid varit så att kommissionen och rådet har arbetat för att förmå de båda förbunden på Cypern att delta i gemensamma projekt .
Det har hittills - som ni vet - inte lyckats , och man har frågat mig om det nu finns några signaler .
Fru Rothe , jag kan uttrycka det så : Jag är övertygad om att ramvillkoren för att uppnå dylika samförstånd har förbättrats väsentligt .
Något accepterande har jag för ögonblicket inte fått .
Det förväntar jag mig inte heller innan vi har gått in i direkta samtal .
Sådana kommer först något senare .
Ramvillkoren har förändrats genom att en hel rad saker som hittills har varit omöjliga nu har gjorts möjliga genom Helsingfors-besluten , men framför allt förstås genom att deltagarnas politiska strategier har genomgått genomgripande förändringar .
Jag har alltid tyckt att den gamla linjen som går ut på att Cypern under alla omständigheter skall upptas först när den politiska konflikten har lösts , att den linjen har en svag punkt , nämligen att den inte är någon övertygande sporre för den turkiska gemenskapen på Cypern att verkligen delta , för enligt denna strategi behövde den turkiska gemenskapen ju inte göra något annat än att luta sig tillbaka och vänta .
Ett medlemskap för Cypern hade då inte blivit aktuellt .
Nu måste de allvarligt räkna med risken att integrerandet av Cypern i Europeiska unionen fullbordas , med de chanser till välstånd och säkerhet som detta för med sig för den grekiska gemenskapen , medan den turkiska gemenskapen , vars välståndsnivå redan ligger mycket lägre , skulle sjunka ännu mer .
Således är det min fasta övertygelse att sporren till att förbinda medlemskapsprocessen med lösningen på konflikten har blivit väldigt mycket starkare efter Helsingfors .
Det är också den idén som har legat bakom .
Fru Rothe , efter dessa få veckor är det fortfarande för tidigt att komma med en utvärdering .
Jag har dock ingen anledning att tro att den nya linjen kommer att misslyckas .
Det finns ingen anledning till det heller .
Inte heller finns det anledning att säga att vi kommer att klara det , men jag kan verkligen säga rent ut att förutsättningarna för att vi skall komma ett steg vidare har förbättrats väsentligt .
En sista punkt : I samtalen med Turkiet spelar Cypernfrågan naturligtvis en roll .
I mitt möte med den turkiska utrikesministern i Bryssel för några veckor sedan bad jag givetvis Turkiet om en positiv och konstruktiv hållning i frågan .
Jag vill bara påpeka en sak : Vi kan inte vara hundraprocentigt säkra - åtminstone är inte jag det - på att man bara behöver trycka på en knapp i Ankara för att allt skall gå vägen på Cypern !
Så enkelt är det verkligen inte , utan vi kommer att bli tvungna att föra intensiva samtal med bägge gemenskaperna för att förmå dem att nå samförstånd .
Det gör vi , kapitalet och programmen för detta finns redan .
Jag behöver - det vill jag bestämt hävda - den budgetförordning som föreligger för beslut för att vi över huvud taget skall kunna sätta igång .
Budgetförordningen är den rättsliga ramen för att ta itu med de prioriteringar som är planerade i partnerskapen för medlemskap för Malta och Cypern .
Så länge vi inte har den kan jag inte dra igång någonting eftersom jag då saknar det rättsliga underlaget .
Om den beklagade bristen på samstämmighet på något sätt skulle ha med denna punkt att göra så måste jag säga att denna förordning bara är en rättslig ram och ingenting annat .
Arbetet med att fylla ut denna rättsliga ram finner ni i prioriteringarna inom partnerskapsavtalen för medlemskap som förra året beslutades av kommission och råd och som nu tillämpas i planeringen och i projektledningen .
Tvärtom skulle jag säga : Det finns många områden inom den europeiska politiken där man kan klaga på bristande samstämmighet .
I detta fall vill jag dock för kommissionens och rådets räkning göra anspråk på att ha utvecklat en mycket tydlig , öppen och samstämmig politik . .
( DE ) Herr talman , herr ordförande !
När nu kommissionären på ett synnerligen samstämmigt vis har förklarat för oss att den bristande samstämmigheten låg hos dåvarande rådsordförande och dennes Europaminister skulle ni kanske kunna hjälpa oss och kommissionären så att detta beslut nu kan fattas .
En lösning som skulle hjälpa vore om ni gav ett positivt svar på min fråga om budgetplanen till 2004 och om rubrik B7 , eller om ni åtminstone ville ge uttryck för att det portugisiska ordförandeskapet avser att anstränga sig för att kompensera den tidigare bristande samstämmigheten - liksom kommissionären kommer att försöka göra i kommissionen . .
( PT ) Herr talman !
Jag tror att den fråga som ställdes av min kollega och gode vän Elmar Brok kommer att övervägas i rådet .
Den kritik som gavs det förra ordförandeskapet är enligt min mening inte relevant .
Jag tror att det som gjordes av det förutvarande ordförandeskapet när det gäller definitionen av budgetplanen var ett utmärkt arbete , oberoende av vem som var involverad i detsamma .
Den fråga som tas upp är i alla fall viktig och vi kommer att fortsätta att ge de förslag som kommissionen lägger fram i den riktningen vårt stöd .
Herr rådsordförande !
Jag har förstått att Brok egentligen menade ett ordförandeskap som ligger ännu längre tillbaka i tiden .
Herr talman !
Jag hade ställt en konkret fråga till Verheugen om finansieringsinstrumentet Meda som han dock inte har svarat på .
Jag vill verkligen be honom att göra det , eftersom även omröstningsförfarandet kring olika ändringsförslag som vi har framför oss beror på hans svar .
Bäste herr Poos , jag ber om ursäkt .
Det fanns en oklarhet just på den punkt som er fråga gällde .
När det gäller Meda är det alltså så att Malta och Cypern kan delta i de överregionala programmen , inte i de landsspecifika eftersom inkomsterna är för höga .
Tack , kommissionär Verheugen !
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum på torsdag .
 
Frågestund ( rådet ) Nästa punkt på föredragningslistan är frågor till rådet ( B5-0009 / 2000 ) .
Fråga nr 1 från ( H-0022 / 00 ) : Angående : Kontroll av oljefartyg som seglar in på gemenskapens vatten Olyckan med oljeutsläppet från tankern Erika orsakade nyligen stora skador längs den franska kusten .
Vilka åtgärder föreslår rådet för att man skall kunna kontrollera oljefartyg som seglar under bekvämlighetsflagg och som inte uppfyller gemenskapens säkerhetsbestämmelser då de seglar in på gemenskapens vatten ?
Herr talman , ärade kollegor !
Den 24 januari snubblade rådet på konsekvenserna efter tankfartyget Erikas förlisning månaden innan .
När rådet i det läget såg hur upprörd allmänheten blev av händelsens förödande konsekvenser uttalade man sin oro vad gäller tankfartygens säkerhet och det miljöskydd som borde förknippas med denna .
Rådet var varken okänslig för den här typen av frågor eller för behovet att vidta kompletterande åtgärder .
Man underströk hur viktigt det var för rådet att vidta nya åtgärder på gemenskapsnivå , men även när det gällde sitt eget arbete tillsammans med de internationella organisationerna .
Som alla vet så ser dagens gemenskapslagstiftning till att hamnmyndigheterna förrättar inspektioner ombord på alla utländska fartyg , inklusive dem som stoltserar med konvenansflagg .
Uppfylls inte de internationella normerna kvarhåller man fartygen .
Det finns ett direktiv som sedan 1995 reglerar detta .
När det gäller framtiden så noterade rådet att funderingarna på kommissionsnivå snart kommer att resultera i ett nytt uttalande om säkerhet för tankfartyg och i nya förslag för bättre kontroll i enlighet med inspektionsmyndigheterna .
Man planerar också att förstärka själva strukturen på de tankfartyg som anlägger gemenskapshamnarna .
De här handlingarna följs upp i rådet ( transport ) och jag kan följaktligen , å rådets vägnar , informera er om att vi kommer att fortsätta att prioritera de förslag som kommissionen med största sannolikhet kommer att lägga fram i den här frågan och som vi menar är grundläggande för miljöskyddet .
Givetvis kommer parlamentet att få yttra sig i det här ärendet eftersom det är underställt medbeslutandeförfarandet .
Det gläder mig att rådet betraktar den här frågan som en anledning till eftertanke .
Rådets ordförande kommer från Portugal , ett land som direkt hotas av en situation som denna .
Om vi tänker funderar för länge , kan det hända att ett oljefartyg under liknande omständigheter går på grund utanför Algarve innan sommaren , förstör den portugisiska turistindustrin i sommar , och med litet tur för havsströmmarna föroreningarna vidare till ön Madeira - för strömmarna går åt det hållet - och då störs även turismen på Kanarieöarna .
Tror inte herr rådsordförande att vi bör sluta fundera och i stället vidta kraftåtgärder i den här frågan , med tanke på att vi redan i dag förfogar över metoder för kontroll av den här typen av oljefartyg på öppet hav ?
Historien om Erika är onekligen en historia som ter sig komisk .
Ett franskägt fartyg med maltesisk bekvämlighetsflagg , hinduisk besättning , sjöcertifikat utfärdat av Italien på Sicilien , som senast inspekterades , jag tror det var i Bulgarien .
Fartyget höll på att sjunkna , kaptenen såg att det höll på att sjunkna och förstod att det inte ens skulle nå fram till närmaste hamn .
Jag anser att sådant inte bör tillåtas .
Det kan leda till enorma skador på ert land , herr ordförande , och även på mitt , Spanien .
Ärade kollega !
Jag kan inte låta bli att dela er oro och jag måste få säga att i ett kustland som ordförandeskapets land så är man givetvis djupt oroad över detta - trots att man inte har några egna tankfartyg .
Vi måste dock följa normerna och de är som de är .
Den normgivande ramen är 1995 års direktiv , ett direktiv som har en samling lagar med viss flexibilitet som eventuellt borde gås igenom på ett mera rigoröst sätt .
I det här området måste vi fungera i samklang med övriga världen , det vill säga vi reagerar efter omständigheterna .
Inför situationens allvar borde vi glädja oss åt att myndigheterna åtminstone har reagerat och börjat reflektera över eventuella lagstiftningsåtgärder .
Kommissionens avsikter i det här fallet är bra , man har för avsikt att förstärka tillämpningen av 1995 års direktiv .
Rådet vill gärna se att den här frågan prioriteras i rådet ( transport ) och vår avsikt är att snabbt behandla den .
Vi hoppas också att frågan lika snabbt kan tas upp i Europaparlamentet genom ett medbeslutandeförfarande .
Herr talman !
I Kotka i Finland ligger för närvarande ett fartyg lastat med kemikalier som seglar under bekvämlighetsflagg .
Fartyget ligger för ankar utanför hamnen eftersom det på grund av det skick som det befinner sig i utgör en säkerhetsrisk för hamnen och närliggande områden och eftersom man i brist på finansiärer inte kan slutföra fartygsinspektionen .
Har EU några som helst möjligheter att skapa ett enhetligt inspektionssystem där man även garanterar betalning från gemenskapens medel för de fartyg under bekvämlighetsflagg som inte själva kan betala ?
Ärade kollega !
Som ni förstår har jag inte den information som behövs för att ge er ett korrekt svar tillgänglig just nu .
Den information som finns tillgänglig har att göra med 1995 års direktiv och där har man inte vidtagit några åtgärder i den riktningen .
Rådet kommer i alla fall att ge er ett konkret svar om de möjligheter som står till buds också gäller för det här fallet .
Fråga nr 2 från ( H-0024 / 00 ) : Angående : Hög barnadödlighet i Kosovo Enligt Världshälsoorganisationens senaste uppgifter till FN har Kosovo högst barnadödlighet i Europa ; nästan 50 procent av alla för tidigt födda barn dör .
Till följd av kriget har missfallen ökat kraftigt och de barn som inte föds för tidigt är mindre utvecklade än normalt .
Kan rådet , mot bakgrund av den humanitära hjälp som EU tillhandahåller och det politiska sändebudet Bernard Koushners ansträngningar , meddela vilka åtgärder det har vidtagit till skydd för kvinnorna i Kosovos rätt till moderskap och för gravida och födande kvinnors samt spädbarns hälsa ?
Herr talman !
Ledamot Karamanous fråga är en fråga av största betydelse vilket vi inte kan bortse från .
Vi är fullständigt medvetna om den svåra och dramatiska situation som människorna i Kosovo befinner sig i och problemet för dem som har förflyttats inom regionen men som härstammar från Kosovo och konsekvenserna av detta när det gäller till exempel barnens hälsa och dödsfrekvensen .
Det är uppenbart att Europeiska unionen klart och tydligt har bistått det internationella samfundets ansträngningar att tillhandahålla humanitärt stöd .
Som ni vet så bidrog Europeiska gemenskapen med totalt 378 miljoner euro bara till provinsen Kosovo , till detta kan man tillägga medlemsländernas egna nationella bidrag .
Bidraget omfattar flera olika projekt inom området för hälsa , som exempelvis vattensaneringen .
Utöver detta ger Europeiska unionen som vi alla vet ett stöd till Förenta nationernas flyktingkommissariat , vilket 1999 uppgick till 66,3 miljoner euro .
Jag tror att ledamoten vet att man på grund av en nödvändig arbetsfördelning mellan de internationella givarna överlämnade hälsosektorn i Kosovo till Världshälsoorganisationen .
Organisationen är fullständigt medveten om den alarmerande situationen när det gäller barns hälsa och man har koncentrerat sina ansträngningar på att förbättra de grundläggande förhållandena på förlossningskliniker och andra sjukhus .
Vi är medvetna om att situationen inte på långa när är löst på ett tillfredsställande sätt , att den är självverkande och har en dimension som förutom barnens hälsa även påverkar andra hälsoområden .
Det är en politisk situation , inte enbart en teknisk , det har att göra med en lösning av den politiska situationen , eftersom det också här finns dimensioner som inte bör förglömmas och som har påverkat det som fram till nu är det internationella samfundets oförmåga att organisera ett multi-etniskt samhälle i Kosovo , vilket fatalt har påverkat hur hälsosystemet har förbättrats i regionen .
Tack , herr rådsordförande , för ert svar , som kompletterar det som kommissionär Patten i går sade i frågan .
Dock har , herr ordförande , den summa på 378 miljoner euro som ni sade att man gav under 1999 i själva verket visat sig vara helt otillräcklig för att skapa grundläggande människovärdiga förhållanden i Kosovo , i synnerhet när det gäller tillhandahållande av hälsotjänster .
Anser ni inte , herr rådsordförande , att bara det faktum att barndödligheten har ökat utgör en skandal för den europeiska kontinenten , en skam , som borde aktivera oss alla , så att den hjälp som vi tillhandahåller blir effektivare och generösare ?
Situationen var naturligtvis inte idyllisk före bombningarna , tvärtom , skulle jag säga , men det skedde en tydlig försämring av både den fysiska och den mänskliga miljön efter Natos attacker .
Är det följaktligen inte , herr rådsordförande , en fråga av moralisk karaktär för oss att försöka skapa människovärdiga förhållanden för de hårt prövade invånarna i Kosovo och , framför allt , att genomföra vad vi har lovat dem ?
Ärade kollega !
Jag erkänner att alla bemödanden som har gjorts i Kosovo har varit otillräckliga .
Jag tror inte att någon av oss tvivlar på detta .
Jag vill inte koppla ihop den här frågan med kommentarerna om perioden " före " och " efter " Natos intervention .
Vi kommer förmodligen att ta upp den frågan vid ett senare tillfälle .
Jag vill dock nämna att vi i Europeiska unionen är medvetna om att vi gjort vad vi kunnat med de finansiella medel som står till vårt förfogande för Kosovo .
Tänk på att vårt ansvar i regionen är ett med det internationella samfundet delat ansvar .
Det är ett ansvar där Europeiska unionen har en särskild uppgift , och vi kan inte göra anspråk på att snabbt bygga upp strukturer som , precis som ledamoten nämnde , redan före det militära ingripandet i Kosovo inte var de bästa .
Ärade kollega , jag tycker inte att de militära aktionerna i Kosovo signifikativt har förstört strukturerna för folkhälsan utan de har mera direkt påverkat den aktuella situationen .
Den aktuella situationen har huvudsakligen att göra med det dramatiska läget för människor på flykt , den har att göra med ekonomiska frågor och hur de grundläggande hälsobehoven tillgodoses efter den globala avregleringen av den organisatoriska administrationen i Kosovo .
Det är primärt detta som ligger till grund för den aktuella situationen .
Så länge vi inte löser den politiska situationen , vilket måste göras genom en resolution av Förenta nationerna , så går inte barnhälsoproblemet att lösa , och det kommer heller inte att finnas någon lösning för andra utvecklingsområden i regionen .
Jag skulle vilja bredda debatten något till situationen i Mitrovica .
Där har världssamfundet , även med europeisk medverkan , återuppbyggt sjukhuset , men det ligger i den norra delen av staden , vilket gör det mycket svårt för kosovoalbaner att få tillträde till detta sjukhus .
Det innebär således att kosovoalbanerna även fortsättningsvis är utstötta från all medicinsk vård .
Det sker också på andra platser i landet , vilket gör att det är spänt mellan kosovoalbaner och serber , att ingen längre litar på någon och att kosovoalbaner inte vill bli vårdade av serber och omvänt .
Jag förstår verkligen att ni säger , och det gör ni med rätta , att Europeiska unionen måste samarbeta i större internationella sammanhang .
Men vad kommer ni att lägga tyngdpunkten på ?
Vad kommer ni att göra för att se till att kosovoalbanerna kan få omvårdnad på ett sjukhus , bland annat i det i Mitrovica ?
Matrovicas fråga känner vi igen , ärade kollega .
Det är fråga om en mycket speciell situation med vissa inter-etniska konflikter som lyckligtvis inte är så allvarliga i andra områden i Kosovo .
Jag har full förståelse för ledamoten .
Jag vill dock nämna att det som Bernard Kouchener har gjort i den här frågan ligger i linje med Förenta nationernas resolution , man har försökt skapa förutsättningar för multi-etniska strukturer som på olika administrativa nivåer kan gagna flera samfund .
Jag tycker inte att vi i den här frågan skall dra förhastade slutsatser om ansvaret , för ansvar har många .
Situationen i Matrovica är beklagansvärd , läget är synnerligen spänt , men jag tror att de åtgärder som i sista stund har vidtagits för att få området säkert är positivt .
Jag vill dock påpeka att vi tyvärr inte kan bistå med någon polisiär styrka - vilket har att göra med medlemsländernas bidrag - för att garantera det som vi föresatte oss att göra med en postmilitär aktion , det vill säga att bygga upp tillräckligt säkra inter-etniska samordningsmekanismer för de olika folkgrupperna så att de får tillträde till sjukhusen .
Fråga nr 3 från ( H-0027 / 00 ) : Angående : Åtal mot Nato i krigsförbrytartribunalen Människorättsorganisationer såsom " Human Rights Watch " i USA har redan samlat in avsevärda uppgifter om brott som Nato begått i samband med bombningarna i Kosovo och Serbien , i syfte att väcka talan i krigsförbrytartribunalen i Haag .
På grundval av dessa uppgifter , som till viss del redan har lagts fram i domstolen , anklagas Nato för allvarliga brott mot internationella mänskliga rättigheter och överlagt mord .
Anser rådet att denna typ av anklagelser bör anföras i krigsförbrytartribunalen för en grundlig rättslig undersökning ?
Om en rättslig undersökning av anklagelserna mot Nato skulle äga rum , hur har rådet då för avsikt att handla i fråga om den höge representanten för GUSP som under krisperioden var Natos generalsekreterare ?
Finns det möjlighet att avstänga honom från sin befattning till det att den rättsliga undersökningen slutförts ? .
( PT ) Herr talman !
Ledamot Alexandros Alavanos fråga väcker funderingar av en mera global karaktär .
Rådet har vid ett flertal tillfällen visat att man var övertygad om att Nato såväl var tvungen som berättigad att vidta de kraftiga åtgärder som vidtogs för att avvärja extremistaktioner , aktioner som klart och tydlig kränker Förenta nationernas säkerhetsråds resolutioner .
Jag förstår att man kan tolka Natos agerande och legitimiteten av detta på olika sätt .
Alla är vi fria att tycka vad vi vill .
I mitt land hade de olika parlamentariska grupperna olika åsikter .
Det är som det är .
För rådet står det i alla fall klart att målet med Nordatlantiska fördragsorganisationens flygräd över Förbundsrepubliken Jugoslavien var att sätta stopp för den humanitära katastrofen i Kosovo förorsakad av regimen i Belgrad .
När rådet ( allmänna frågor ) i Luxemburg godkände ståndpunkten den 8 april åskådliggjordes målet klart och tydligt .
Natos åtgärder vidtogs inte med glädje , vilket måste framgå , och de genomfördes bara som en sista utväg när det var uppenbart att alla möjligheter till en fredlig lösning var uttömda och myndigheterna i Belgrad höll på att samla sina styrkor för att driva bort kosovoalbanerna från sitt territorium .
Ledamoten vet säkert att åklagaren vid sitt senaste besök på Natos högkvarter påpekade att den internationella domstolen är tvungen att granska alla anklagelser , inklusive dem som har formulerats mot Nato av kanadensiska fredsgrupper .
En sådan obligatorisk granskning skulle genomföras allteftersom anklagelserna gjordes .
Jag har i alla fall med mig ett uttalande av åklagaren där hon säger att Natos aktioner inte är underställda någon granskning av åklagaren vid den internationella brottmålsdomstolen för före detta Jugoslavien , och att det inte finns någon formell granskning av Natos aktioner i Kosovokonflikten .
All information som mottagits under de senaste sex månaderna , må vara av privatpersoner eller av grupper som begär att Natos aktiviteter under Kososvokonflikten granskas , registrerades av åklagaren .
Informationen kommer givetvis att analyseras av åklagaren och tids nog får vi veta om det finns skäl att agera eller inte .
Åklagaren har hittills valt att inte behandla anklagelserna mot Nato .
Jag tackar rådsordföranden , men jag håller inte med honom om att Natos ingripande var avsett att stoppa en humanitär katastrof , för vi har även i dag en humanitär katastrof i Kosovo , och Milosevic inferno följdes av UCK : s och Natostyrkornas inferno .
Och kanske har även rådsordföranden noterat att nära hälften av de frågor som han skall svara på i dag handlar om Kosovo .
Icke desto mindre håller även rådsordföranden med om att frågan om en undersökningsprocess mot Nato i krigsförbrytardomstolen , efter en anmälan från bland annat kanadensiska fredsorganisationer , är öppen .
Och min fråga , på vilken rådsordföranden inte gav något svar , är följande : Om denna undersökningsprocess inleds , i vilken den huvudsaklige eller , om ni vill , en av de huvudsakliga undersökta - och troligtvis skyldiga - kommer att vara Solana , som i dag är " hög representant för Europeiska unionens gemensamma utrikes- och säkerhetspolitik " , borde i så fall inte , om detta inträffar - och domstolens allmänna åklagare är positiv till att starta processen - , borde då inte Solanas befogenheter suspenderas , åtminstone till dess att hans oskuld är bevisad ?
Ärade kollega !
I händelse av att man försöker agera på det här sättet mot Nato och i fall en sådan händelse skulle personifieras i Javier Solana , så måste vi vara medvetna om att Javier Solana innehar ett annat ämbete i dag .
Det ämbete han i dag innehar har absolut inget att göra med det tjänsteåligganden han då hade som Natos generalsekreterare .
Finns det ingen internationell domstolsmyndighet som på något sätt kan rättfärdiga definitionen av brott genom angivandet av Javier Solana , något som inte har inträffat på långa vägar , så kommer givetvis Europeiska unionen inte att inta någon som helst ståndpunkt i den här frågan .
Herr talman !
Jag tror att Alavanos förväxlar Nato och Milosevic .
Milosevic borde ställas inför krigsförbrytartribunalen , och Nato borde vi ge Sacharovpriset !
Men jag har en helt annan fråga till rådet .
Hur ser det ut med uppbyggnaden av förvaltning och rättsväsende och framför allt polisen i Kosovo ?
Ni antydde det nyss , här står vi inför en katastrof , och ingenting görs .
Här måste planeras ett raskt agerande !
Jag vill först och främst säga att jag instämmer med ledamoten när det gäller att prioritera identifieringen av personer som kan ställas till svars .
När det gäller den juridiska uppbyggnaden av Kosovo så har vi ett flertal gånger haft tillfälle att höra Bernard Kouchners beskrivning av hur svårt det är att bygga upp ett administrativt maskineri och en rättslig struktur .
Vi vet att de första stegen togs för flera månader sedan .
Svårigheterna känner vi till , särskilt de finansiella .
De svårigheter som Bernard Kouchner har stött på vid den administrativa uppbyggnaden känner vi också till , i synnerhet svårigheterna med att rekrytera polisstyrkor för den dagliga säkerheten .
Ärade kollega , det är ett ansvar som vi måste ta och fundera över inom Europeiska unionen .
I måndags i rådet ( allmänna frågor ) togs Kosovofrågan upp ett antal gånger .
Efter en del uttalanden utövades påtryckningar på de medlemsländer som hade lovat att ställa upp med polisiära styrkor men inte fullgjort sina åtaganden .
Några av medlemsländerna försökte ursäkta sig med att de redan har militära styrkor på plats och att man inte hade kunnat komplettera med de polisiära styrkorna så snabbt som man hade velat .
Jag är fortfarande övertygad om att detta kommer att vara det som på ett avgörande sätt kommer att misskreditera Bernard Kouchners arbete samt regleringen och normaliseringen av den administrativa strukturen i Kosovo , i synnerhet den rätttsliga och polisiära .
Detta kommer att ha fatala konsekvenser , klara och tydliga när det gäller vår förmåga att reglera den inter-etniska samordningen .
Vi vet alla att om inga åtgärder vidtas inom kort kommer konflikter att uppstå , precis som de vi såg för några timmar sedan och de kommer att spridas till andra områden i Kosovo .
Det här är en fråga som i första hand berör Nato , men som Europeiska unionen inte har svårt att ansluta sig till eftersom man delar Natos uppfattning i de här frågorna .
Jag vill att detta skall stå klart , det är rådets ståndpunkt och det bör inte råda några tvivel om detta .
Ledamoten är medveten om hur svårt det är att först och främst välja mål vid en militärinsats , i synnerhet när det gäller flyganfall .
Han är också medveten om att det finns mål som inte är militära mål utan infrastrukturella mål , vars syfte är att förekomma militärstyrkornas verksamhet .
Här kommer vi uppenbart in på ett område , ett grått område , där ledamoten kommer att säga att civila mål är mål som exempelvis broar , väg- och järnvägsnät medan andra säger att detta är militära mål , eftersom de bistår de militära strukturerna vid aggressiva insatser , insatser som de som Milosevics styrkor genomförde i Kosovo .
Vi tolkar detta på olika sätt , det är några mål som skiljer oss åt .
Tyvärr var det också så som alla tolkade militärinsatserna i Kosovo .
Det fanns vissa civila sektorer , sektorer som hade att göra med infrastruktur med direkt anknytning till folket och det fanns till och med befolkade områden som träffades under Natos lufträder .
Vi vet , det inträffar i alla krig och kriget i Kosovo är inte ett rent krig , ett föredömligt krig , det är ett möjligt krig .
Det var bara det att det var ett nödvändigt krig .
Förutom att det var ett möjligt krig , var det nödvändigt för att sätta stopp för en absolut oacceptabel aggression avskydd av hela det internationella samfundet .
Ärade kollega , oavsett vilken tolkning vi gör i efterhand - görs inget så är det lätt att göra tolkningar i efterhand - så tror jag att om man tittar på det som hände i Bosnien-Herzegovina och på den strafflöshet och förlängningen av denna som situationen i Bosnien-Herzegovina förorsakade , så kan vi kanske se Natos militära insats i Kosovo som litet mindre ödesdiger .
Fråga nr 4 från ( H-0028 / 00 ) : Angående : Den turkiska blockaden av Armenien När nu en gång Europeiska unionen med hjälp av det partnerskaps- och samarbetsavtal med Armenien som undertecknades den 12 oktober 1999 aktivt verkar till förmån för sociala , ekonomiska och politiska relationer med Armenien , vad gör rådet för att söka förmå Turkiets regering att upphäva den ekonomiska blockaden av Armenien ?
Är det dags för Turkiets regering att att upphäva den ekonomiska blockaden av Armenien ? .
( PT ) Herr talman !
Anledningen till ledamotens fråga är en regional konflikt , om man läser mellan raderna , samt förmodandet att det finns en bilateral förbindelse som har att göra med Armenien och Turkiet .
Det som ligger bakom den här frågan är uppenbart frågan om Nagorno Karabach samt konflikten mellan Armenien och Azerbajdzjan , som tack vare de goda förbindelserna mellan Azerbajdzjan och Turkiet givetvis har sina konsekvenser .
Apropå den här förbindelsen mellan Europeiska unionen och Armenien , eftersom det är den som kan intressera oss , så vill jag säga att ikraftträdandet av avtalet om intresseföreningar och samarbete i juli 1999 och det första sammanträdet i oktober i fjol visar hur pass viktiga förbindelserna med Armenien är för Europeiska unionen .
Ett av målen är utvidgandet av handelsförbindelserna , i synnerhet när det gäller handel och investeringar samt möjligheten att hålla en bilateral politisk dialog med Armenien då landet spelar en viktig roll i regionen .
Som sagt , frågan om Nagorno Karabach är fortfarande en fråga som är viktig att lösa och som naturligtvis försvårar stabiliteten i södra Kaukasus .
Som första prioritet måste vi enligt vår mening intensifiera alla åtgärder så att konflikten kan lösas .
Europeiska unionen har vidtagit åtgärder för att underlätta processen och givetvis är vi medvetna om att också Turkiet måste vara konstruktiv i den här frågan och ta på sig ett stort ansvar .
Turkiet togs i december 1999 upp som kandidatland till Europeiska unionen .
Den politiska dialogen med Turkiet kommer att intensifieras i och med den nya situationen .
Som företrädare för Europeiska unionens ordförandeskap var jag i Ankara i anslutning till beslutet och det meddelande vi lämnade de turkiska myndigheterna var att den politiska dialogen är av synnerligen stor vikt och att vi vill dra nytta av Turkiets roll i regionen , i synnerhet när det gäller förbindelserna med Centralasien och Kaukasus .
Inom ramen för de här förbindelserna med Turkiet som vi gärna ser politiskt privilegieras , främst tack vare landets position i regionen och det viktiga geostrategiska läget , måste vi försöka nå samstämmighet i de internationella frågorna .
Vi förväntar oss att Turkiet intar en konstruktiv attityd , en positiv attityd .
Vi hoppas särskilt att Turkiet , inom ramen för den politiska dialog som föregår det förfarande som kan leda fram till förhandlingarnas början , kan ansluta sig till Europeiska unionens uttalande om den gemensamma utrikes- och säkerhetspolitiken .
Här är jag övertygad om att Turkiet inte kan undvika den tolkning vi har gjort om nödvändigheten av att finna rimliga lösningar för Nagorno Karabach , lösningar som beaktar såväl de lagliga aspekterna för Armenien som för Azerbajdzjan .
Herr talman !
Jag vill tacka företrädaren för ordförandeskapet för hans svar .
Dock är jag ledsen att man visserligen i första hand ser detta bilateralt men att det till slut ändå är ett triangelförhållande .
Vi beviljar partnerskapsbidrag och har samarbetsavtal för att hjälpa Armenien , och trots det kan ju hjälpen inte alls bli effektiv eftersom Turkiet genomför en handelsblockad , så att armenierna på många punkter över huvudtaget inte kan komma framåt .
Med Turkiet förhandlas det om ett eventuellt medlemskap , och det ligger ju i allas vårt intresse att varje stat som vill bli medlem också vårdar fredliga förbindelser med sina grannar längs gränserna .
Kan ni inte öka trycket på Turkiet för att möjliggöra en fredlig utveckling , för att också ge armenierna en chans till den utveckling som är nödvändig för att samarbetet skall kunna gå vidare ?
Ledamoten har rätt när hon säger att vi måste använda förbindelserna med Turkiet just för att få landet att agera konstruktivt , i synnerhet när landet blir en del av lösningen och inte en del av problemet .
Tack vare att Turkiet har gått in i en ny fas i sina förbindelser med Europeiska unionen och tack vare att Turkiet nu måste konfronteras med Europeiska unionens ställningstagande i den gemensamma utrikes- och säkerhetspolitiken så tror vi , och det här kan vi inte dölja , att vi på det här viset kan testa Turkiets inställning till Europeiska unionens utrikespolitiska prioriteringar .
Givetvis är förbindelserna med Armenien , som fjolårets avtal är ett bevis på , en del av den utrikespolitiken .
Vill Turkiet dela Europeiska unionens grundläggande värderingar och unionens allmänna förbindelseramar - oberoende av den bilaterala idiosynkrasi man eventuellt kan ha inför ett annat land , så måste Turkiet generellt sett följa de grundläggande ramarna för Europeiska unionens utrikesförbindelser .
Vi är övertygade om att man mycket snart kommer att prioritera den här frågan i de bilaterala förbindelserna mellan Europeiska unionen och Turkiet .
Eftersom de behandlar samma ämne , kommer frågorna 5 och 6 att tas upp tillsammans : Fråga nr 5 från ( H-0031 / 00 ) : Angående : Förvärrad situation i Kosovo Folkmordet på serber och andra icke-albanska , etniska grupper i Kosovo har förvärrats .
Till och med Bernard Koushner tillkännagav nyligen att den politiska situationen och säkerhetsförhållandena i området inte alls är tillfredsställande .
Det har också uttryckts klagomål över att FN : s resolution nr 1244 inte har efterlevts .
Resolutionens föreskrifter om garantier för alla invånare i Kosovo har inte följts , extremistiska utbrytarstyrkor främjas och som kulmen på problemen har den förre UCK-ledaren H. Thaci utnämnts till tillförordnad premiärminister för Kosovo och UCK till Kosovos skyddsstyrka .
Vilka åtgärder har rådet mot bakgrund av ovanstående för avsikt att vidta för att FN : s beslut , i synnerhet resolution nr 1244 , skall efterlevas och för att förhindra att provinsen Kosovo bryter sig ur Serbien ?
Fråga nr 6 från ( H-0122 / 00 ) : Angående : Etnisk rensning av serber i Kosovo Natos och EU : s bombningar av Jugoslavien motiverades med att man ville sätta stopp för den etniska rensning av kosovoalbaner som Serbien hade gjort sig skyldigt till .
Sedan dessa bombningar upphörde , och sedan Kfor-styrkan upprättades den 12 juni 1999 , har 200 000 serber bosatta i Kosovo fördrivits och 768 mördats .
Sålunda har rensningen av serber varit jämförelsevis större än rensningen av kosovoalbaner .
Under de senaste dagarna har vi sett hur serber mördas av kosovoalbanska maffior utan att dessa gärningar bestraffas på något sätt .
Vilket beslut ämnar rådet fatta för att en gång för all sätta stopp för denna form av etnisk rensning och för att garantera respekt för mänskliga rättigheter för samtliga befolkningsgrupper i Kosovo , oberoende av etniskt ursprung eller religion ?
Herr talman !
Som jag tidigare tog upp så är situationen i Kosovo ett problem som man i måndags uppmärksammade i rådet ( allmänna frågor ) .
Rådet sade sig stödja Unemic och generalsekreterarens sändebud , Bernard Kouchner , i arbetet med att inrätta en interimsadministration i Kosovo och där man garanterar att alla styrkor skall vara inkluderade , framför allt de som hittills har vägrat att vara en del av denna interimsstruktur .
Den höga representanten för den gemensamma utrikes- och säkerhetspolitiken , Javier Solana , visade ministerrådet för allmänna frågor en utvärdering av situationen och efter denna inväntas nu förslag , i synnerhet förslag på åtgärder för en intern justering som inte bara skall tillåta en viss flexibilitet i de interetniska förbindelserna utan också - som jag redan tidigare nämnde - ett inrättande av nya polisiära strukturer och system så att situationen i Kosovo inte skall förvärras när det gäller maktmissbruk , narkotikahandel och kriminalitet , något som den nuvarande styrkan inte har lyckats med .
Ärade kollega , därför är ministerrådet synnerligen oroad över den aktuella situationen i Kosovo .
Man är särskilt oroad över den serbiska befolkningens massutvandring och över andra etniska och religiösa minoritetsgruppers situation ( minoriteter som många gånger inte nämns tillräckligt mycket när man talar om diskrimineringen i Kosovo ) .
Man är också besviken och oroad över det interetniska våldet som man fortfarande kan notera .
Som jag tidigare fick tillfälle att säga så är den nya antagonismen i Mitrovica bara ett exempel på de svårigheter som måste övervinnas när det gäller det under årtionden ackumulerade misstroendet .
Vi befinner oss just nu bara i en fas i en process med flera faser i förfluten tid , och jag tror att vi alltid måste titta på den i ett historiskt perspektiv .
Europeiska rådet visade otaliga gånger att man ville skapa ett demokratiskt och multietniskt Kosovo i enlighet med resolution 12 / 44 av Förenta nationernas säkerhetsråd .
I synnerhet vill man se att alla flyktingar säkert och utan hinder kan återvända .
Ärade kollega , för oss är detta fortfarande en central fråga för vårt engagemang i regionen , oavsett de tvivel som resolution 12 / 44 kan ha väckt , och låt detta stå klart .
När det gäller det som är till skada för regionen så vill jag säga att rådet fördömer alla våldsgärningar , all förföljelse och intolerans oavsett gärningsman .
Som svar på den aktuella situationen stöder rådet till fullo Förenta nationernas uppdrag i Kosovo .
UNMIK står för de budgeterade medlen och för den så kallade " UNMIK : s fjärde pelare " , som har att göra med återuppbyggnaden och den ekonomiska rehabiliteringen .
För att utvärdera de framsteg som hittills gjorts av UNMIK måste man komma ihåg att den situation man befinner sig i är extremt svår , det vill säga en stor mängd flyktingar och omplacerade måste få komma tillbaks , en nästan totalförstörd infrastruktur , en radikalisering som fortfarande är mycket aktiv inom alla sektorer i Kosovo , en ekonomisk kollaps , en total frånvaro av interna inkomster och administrativa strukturer på lokal- och distriktsnivå vilka helt har brutit samman , liksom rätts- och polisväsendet .
Boven i dramat är kriget och ett årtionde av försumlighet efter Belgrads avskaffande av Kosovos självstyre .
Detta är viktigt , vi måste komma ihåg att det var Kosovos ändrade författning inom ramen för Republiken Jugoslavien som var orsak till att de etniska konflikterna ökade och ledde till den nuvarande situationen .
Det här får vi inte glömma bort , så att inte tidigare händelser glöms bort av ansvariga historiker .
Under sådana omständigheter menar jag att UNMIK tillsammans med andra inblandade myndigheter och internationella organisationer har gjort vissa framsteg beträffande de mål som nämns i resolution 12 / 44 , även om vi har långt kvar till en tillfredsställande lösning av situationen .
Rådet stöder ändå det särskilda sändebudet Bernard Kouchners beslut att inrätta - som nämnts - ett gemensamt provisoriskt administrativt råd för alla etniska grupper i Kosovo .
Europeiska unionen har försökt få serberna i Kosovo att överväga bojkotten mot nämnda strukturinsats så att ett multietniskt område kan bildas och så att man tillförsäkrar sig en egen plats i den förekommande administrativa strukturen .
Eftersom målet är att bekämpa de multietniska våldet och skapa den säkra miljö som behövs för att förhindra att kosovaner som inte är av albanskt ursprung lämnar provinsen , så stöder å andra sida Europeiska unionen UNMIK : s arbete med att bygga upp en civil polisstyrka av kosovaner .
Trots att bidraget har varit substantiellt måste vi tillstå att Europeiska unionens medlemsländer hittills , som sagt , inte har lyckats utse några konstaplar för nämnda polisstyrka , vilket i högsta grad har inverkat negativt på allmänhetens säkerhet .
Som sagt , i enlighet med de slutsatser som presenterades av rådet ( allmänna frågor ) den 24 januari gör medlemsländerna en kraftansträngning för att finna och komplettera den polisiära styrkan , en ståndpunkt som förnyades av det senaste rådsmötet ( allmänna frågor ) .
En förstärkning av de polisiära styrkorna är också en viktigt uppgift på grund av det ökade hotet från den organiserade brottsligheten .
Kommissionen tänker inkludera kampen mot den organiserade brottsligheten i sitt biståndsprogram för Kosovo år 2000 och man uppmanar medlemsländerna att identifiera vilket typ av bistånd man kan ge för detta .
Vi tror också att en lösning på Kosovos problem - och det är ingen mening att tvivla på detta heller - till stor del är avhängig instabiliteten i de länder som är involverade .
Utan stabilitet kan man inte göra anspråk på att lösa Kosovofrågan .
Lyckas man inte stabilisera den politiska situationen i Albanien - förslag har lagts fram om att kommissionen skall utvärdera hypotesen av ett stabiliserings- och associeringsavtal med Albanien - lyckas man inte stabilisera den politiska situationen i Makedonien i den forna Republiken Jugoslavien och lyckas man inte skapa integrerade modeller för andra områden i det forna Jugoslavien så kommer man inte att klara av att ge Kosovo autonomi .
Det är det globala sammanhanget i regionen och det globala sammanhanget i tillämpningen av stabilitetspakten som kan lösa Kosovos problem .
Herr talman !
Ni får ursäkta mig , men när man lyssnar på rådets företrädare måste man faktiskt fråga sig hur långt skenheligheten , toleransen och delaktigheten kan gå .
Det är ett faktum att man i den hängdes hus , som vi säger i mitt hemland , inte talar om rep .
Jugoslavien var ett fredligt land , en stabilitets- och fredsfaktor .
Med Natos , och i början även Tysklands , attacker blev det som det blev .
Den skyldige är följaktligen inte regeringen i Belgrad , herr talman , utan Nato , imperialisterna med sina attacker .
Hur ser situationen ut i dag ?
Vi har en grov kränkning av säkerhetsrådets resolution 1244 , vilket bevisar att den var en fälla .
350 000 serber , zigenare och andra etniska grupper - dock inga kosovoalbaner - har fördrivits .
900 har mördats , 800 har förts bort med våld ; åtta månader efteråt fortsätter den grova kränkningen av säkerhetsrådets resolution .
Till exempel räcker det inte med att UCK inte avväpnades inom en tremånadersperiod , vilket föreskrevs i resolutionen , utan organisationen har också stick i stäv med Kouchers försäkranden inför Europaparlamentet försetts med modern utrustning och utropats till " Kosovos skyddskår " .
Och jag skulle för att avsluta , herr talman , vilja säga , med anledning av att ministern nämnde Kouchner , att Kouchner med sina 25 påbud kränker Jugoslaviens suveränitet och säkerhetsrådets resolution .
Han har skapat en särskild valuta , en domarkår ...
( Talmannen avbröt talaren . )
Vi måste se verkligheten som den är , herr talman !
Jag tycker inte att ledamoten uttryckte några frågor , han uttryckte några sanningar .
Den första av dem , och som jag noterar här i kammaren , är att Belgrad inte kan ställas till svars för situationen i Kosovo .
Jag ser gärna att detta klargörs för uttalandet är viktigt och av vilket man kan dra slutsatsen att Natos imperialistiska aktiviteter är ansvarig för situationen i Kosovo .
En sällsam tolkning - fast kanske inte alltför sällsam för den delas av de serbiska myndigheterna - men jag tror nog att ledamoten är medveten om att det finns andra tolkningar , och att det internationella samfundet och Europeiska unionens ministerråd har en annan tolkning .
Ärade kollega , om resolution 12 / 44 är en fälla så förstår inte jag heller hur det kan komma sig att ni sedan anser att allt våld i fällan också är negativt .
Resolution 12 / 44 är kanske inte perfekt , men det var den resolution som man kunde enas om för att sätta stopp för en viss bestämd situation .
En resolution som förmodligen fick problem med tillämpningen just av den anledningen att det innebär stabilitet som varken Milosevic eller hans regim har bidragit till .
Jag erkänner , och det gör vi alla , att beteendet hos en del kosovoalbanska styrkor inte heller har varit det bästa och mest intelligenta .
Jag är säker på att Bernard Kouchner på ett konkret sätt även har tagit upp detta .
Vi får inte tro , ärade kollega , att skulden bara ligger på ena sidan och vi får inte tro att vi får glömma det som hänt när vi står i begrepp att analysera rådande situationer .
Sådana här situationer , i synnerhet de på Balkan - ledamoten känner bättre till det här än jag - har alla att göra med det förflutna och med en ackumulering av historiska händelser .
Det finns inte bara " de goda i filmer " .
Situationer av det här slaget är mycket klara - tycker jag - och vi måste alla stå för konsekvenserna och ta på oss ansvaret för vår tidigare tystnad när det gäller Milosevics uppträdande under den tid som han ostraffat kunde göra vad han gjorde , i synnerhet från det ögonblick han återtog självstyret .
( Applåder ) Jag vill tacka för ministerns svar , men samtidigt påminna om att våldet i Kosovo statistiskt sett är större nu än det var före Natos bombningar .
Det är oroväckande att bombningarna har förvärrat situationen , och det bör medges att Nato och Europeiska unionen har agerat felaktigt i och med den åtgärden .
Ministern har talat , och det har han alldeles rätt i - jag håller med om det - om Belgrads skuld i det hela , men man bör också tänka på att underrättelsetjänsten i USA , Tyskland , Frankrike , Italien och Storbritannien har försett UCK , en maffia , med vapen och pengar , och på det viset bidragit till problemen i området .
Därför bär vi alla skulden .
Jag vill ställa en tilläggsfråga på grund av frågans globala natur .
Tror ni inte att det skulle vara en fördel att häva blockaden mot Serbien , så att ekonomin i området normaliserades och att även Kosovo , som en provins i Serbien , skulle ha nytta av det ?
Ärade kollega !
Jag vill bara säga att det är svårt att basera sig på antaganden och sedan uttala sig om vad som hänt om något inte hade hänt .
Varken ledamoten eller jag kan säga vad som skulle ha kunnat inträffa i Kosovo om Nato inte hade bombat .
Och om inte Milosevic och hans regerings allt aggressivare aktioner inte hade lett till en mycket allvarligare situation än den som vi i dag har i Kosovo ...
När det gäller ett lyftande av sanktionerna menar vi , ärade kollega , att Europeiska unionens inställning till Jugoslavien är baserad på en gradvis utvärdering av varje situation .
Vi har satt igång ett energiprogram för att främja demokratin genom att gynna och stödja de kommuner i Jugoslavien som styrs av demokratiska krafter .
I rådet ( allmänna frågor ) reagerade man positivt på den begäran som framställdes av de demokratiska krafterna i Serbien för att för såväl internationella som jugoslaviska flygbolag lyfta embargot .
Detta är ett tecken på Europeiska unionens goda vilja när det gäller situationen i Serbien .
Vi måste förstå att det inte är fråga om att ge de serbiska myndigheterna några förmåner och att det inte är fråga om att ge utan att få något i gengäld .
Såväl de interna mänskliga rättigheterna som det interna politiska systemets funktion i Serbien är under all kritik - och jag hoppas att ledamoten håller med mig om den demokratiska situationen i landet .
Vi ger tillräckligt till Serbien , såväl när det gäller förmåner som lyftandet av sanktioner , dock under förutsättning att Serbien på det internationella planet och i förbindelserna med sina grannländer eller internt uppträder på ett sätt som vi menar följer de grundläggande principerna för det internationella samfundets och de " goda ländernas " uppträdande på det internationella planet .
Herr talman !
Jag är ingen vän till Milosevic eller hans regering .
Icke desto mindre hyser jag de allvarligaste tvivel om legitimiteten för Natos attacker mot Jugoslavien i Kosovo , både med avseende på bristen på bemyndigande från FN : s säkerhetsråd och på grund av att de kunde ha undvikits genom att inte ålägga oacceptabla villkor för Serbiens suveränitet vid Rambouillet .
Den nuvarande situationen i Kosovo , som nu är etiskt rensat på serber och romer , talar för sig själv .
Borde inte Nato åtminstone erkänna skulden för den avsiktliga bombningen av Belgrads TV-torn , vid vilken över 20 civila journalister miste livet , som förblir en stor moralisk skamfläck från kriget och som nu öppnar upp för ett generande eventuellt åtal om krigsförbrytelser mot våra ledare i väst ?
Ärade kollega !
När det gäller Europeiska unionens ståndpunkter så gör man ingen tolkning , ingen selektiv analys av militära mål , som till exempel anfallen mot den infrastruktur som Milosevics politiska system och propaganda kunde stödja sig på .
Därför kan jag följaktligen inte uttala mig om den konkreta situationen och om vi kom överens med Nato eller inte om att utföra den .
Det var en del i en global plan där vi alla var överens .
Några av aktionerna var diskutabla , några erkände Nato själv var beklagliga och andra var av taktiska skäl berättigade för att stoppa Milosevics interna propagandakampanj .
Å rådets vägnar tänker jag i alla fall inte uttala mig om någon specifik militäraktion utförd av Nato .
Herr rådsordförande !
Eftersom jag känner till Balkans historia , skulle jag vilja påminna er om att Jugoslaviens folk under många decennier levde fredligt ihop .
Destabiliseringen började för omkring tio år sedan , i och med Jugoslaviens upplösning , i vilken Europeiska unionen spelade en avgörande roll .
Jugoslaviens brott var att det var det enda landet på Balkan som inte sökte medlemskap i vare sig Nato eller Europeiska unionen .
Vad som nu står kvar efter flygbombningarna , förstörs av det inte alls avväpnade UCK , framför näsan på KFOR , vars roll som ockupationsmakt blir allt tydligare .
Dagligen kommer nya brott mot icke-albanska grupper , men även mot Kosovos kulturella arv , fram i ljuset , liksom hundratals överträdelser av FN : s resolution 1244 .
Enligt min åsikt är det bästa som rådet skulle kunna göra att avbryta ockupationen av denna del av Jugoslavien och söka en lösning som är godtagbar för alla sidor , med respekt för regionens etniska särdrag och - framför allt - med respekt för principen om att man inte blandar sig i andra självständiga länders inre angelägenheter .
Jag har full respekt för ledamotens kännedom och tolkning av situationen i balkan , även om jag har svårt att förstå hur man genom att respektera regionens särdrag kan åstadkomma politisk stabilitet och därmed en lösning på problemet , för om vi tittar på den demokratiska stabiliteten i regionen skulle man kunna säga att det var Jugoslaviens ödeläggelse som orsakade den nuvarande situationen .
Låt oss inte försöka oss på att tolka en internationell manöver .
Jag vill påstå att Jugoslavien var vad det var , en stat med en viss förenlighet i den etniska differentieringen , en stat med en politisk inramning som ur en demokratisk synvinkel var allt annat än idealisk , något som måste stå klart för alla .
Delningen av Jugoslavien är förmodligen ett historiskt faktum som vi måste lära oss att leva med , oavsett begångna misstag litet här och där .
Vi tror inte alls att en reträtt av de internationella styrkorna just nu skulle vara en lösning .
Tvärtom skulle den vara till skada .
Herr talman !
Jag blev litet besviken över det svar som rådsordföranden gav min kollega .
Det är mycket viktigt , om vi betonar att Europa skall vara ett värderingarnas Europa , att vi inte börjar påstå att medlen helgar ändamålen .
Om civila mål bombades och förstördes - att döda civila är olagligt enligt alla mått mätt .
Det bör inte försvaras ens av de av oss som djupt beklagar Milosevicregimen .
Detta är dock inte min fråga .
Min fråga handlar om politiska fångar som hålls fångna i Serbien nu .
Det finns , tror jag , för närvarande omkring 5 000 kosovanska politiska fångar som hålls fångna i Serbien .
Min fråga till rådsordförande är följande .
För det första , är rådet fullt medvetet om och intresserat av dessa fångars öde ?
För det andra , vad har det för avsikt att göra för dem ?
Ärade kollega !
Jag vill börja med att kommentera det jag sade tidigare .
Jag försvarade inte alls anfallen mot civilbefolkningen .
Det jag sade och det jag redan har förklarat är att det finns civila mål som har att göra med strukturer som är en del av den militära aktionen , och ledamoten vet lika väl som jag att en del militäraktioner inte bara riktas mot militära mål , de riktar sig också mot civila mål som komplement till de militära .
Det är uppenbart att vi befinner oss i en gråzon när det gäller vad som är och inte är legitima mål .
Som sagt , låt oss inte bedöma specifika aktioner .
Vi gör en global bedömning av Natos aktioner och den globala bedömningen är positiv och vi delar Natos uppfattning .
När det gäller de politiska fångarna i Serbien , ärade kollega , så är det uppenbart att när jag talar om Serbien av i dag så följer inte Milosevic på det internationella planet de regler som gäller i ett anständigt samhälle .
Jag tänker på Milosevics förhållande till sina medborgare , men framför allt hans sätt att hantera de politiska fångarna , de demokratiska kränkningarna , kränkningarna mot rätten till oppositionell massmedia , kränkningarna mot rätten för icke-statliga organisationer att agera och främja de mänskliga rättigheterna .
Detta är trots allt bara en aspekt av Milosevics skadliga agerande i det jugoslaviska samhället och Europeiska unionen är givetvis bekymrad över situationen .
Därför vill Europeiska unionen fortsätta med sina sanktioner så länge som Jugoslavien internationellt sett inte ändrar sitt uppförande och börjar respektera de värderingar som vi anser vara betydelsefulla .
Fråga nr 7 från ( H-0035 / 00 ) : Angående : Utkastet till en stadga om grundläggande rättigheter Det civila samhället ser med tillfredsställelse på utkastet till en stadga om grundläggande rättigheter och förhoppningen är att denna skall kunna anta de utmaningar som Europa kommer att ställas inför under det 21 : a århundradet .
Kan rådet mot denna bakgrund svara på följande frågor : Hur ser rådet på innehållet i stadgan ?
Vem skall stadgan gälla ?
Medborgare i Europeiska unionen eller i alla europeiska länder , med tanke på utvidgningen ?
Kommer den även att omfatta invandrare o.s.v. ?
Kommer stadgan att befästa Europeiska unionens sociala rättigheter eller kommer den att ha en bredare karaktär ?
Vilka mekanismer kommer att användas i stadgan för att tydligt säkerställa jämlikhet mellan de båda könen ?
Vad anser rådet om att införa stadgan i EU-fördraget ? .
( PT ) Dokumentet om de grundläggande friheterna är en av de viktigare frågor vi arbetar med på institutionsnivå inom Europeiska unionen .
Som ni vet har dokumentet sitt ursprung i det beslut som togs i Köln av Europeiska rådet .
Vi menar att dokumentet är grundläggande för att skapa det som kan betraktas som Europeiska unionens etiska pelare och det som kan betraktas som ett behov för Europeiska unionen på vägen mot en union med värderingar , för att kunna förstärka dimensionen , inte bara internt utan till och med för att legitimera sitt eget externa bejakande baserat på gemensamma värderingar .
Detta är givetvis av stor vikt för de femton .
För fyra , fem månader sedan trodde vi inte att det skulle vara så viktigt för unionen .
I dag tänker vi tack och lov på ett annat sätt , åtminstone några av oss .
Det kommer också att vara betydelsefullt för en utvidgad union , i synnerhet för den framtida kulturpolitiken .
Beträffande dokumentets innehåll : Som ni vet så håller vi fortfarande på att diskutera stadgan .
Två sammanträden har hållits av den grupp som har till uppdrag att utforma den , en grupp som nu kallas konventet för Europeiska unionens stadga för de mänskliga rättigheterna .
Ett flertal problem har dykt upp .
Först och främst måste vi veta om texten är förklarande eller om texten är bindande .
För det andra , stadgans innehåll : oavsett om stadgan är bindande eller inte så har vi ändå ett innehållsmässigt problem , det vill säga om det handlar om en kumulation av ett antal principer som unionens medlemsstater tar i försvar och som finns medtagna i deras interna författningar eller om det är fråga om en ny korpus som på något sätt kan vara unionens gemensamma grundtanke .
Sedan har vi ett annat grundläggande problem , som för övrigt finns med i frågeställningen och som jag tycker är av stor vikt , men som ännu är olöst .
Vi måste ta reda på om stadgan skall tillämpas på unionens medborgare eller om det skall tillämpas på tredje lands medborgare bosatta inom unionen .
Det är också en fråga som ligger på bordet .
Till sist har vi också ett mera svårlöst problem , frågan om rättsordningarnas underställelse , frågan om förenlighet mellan Strasbourgdomstolens rättsordning och Luxemburgdomstolens rättsordning .
Ett problem som måste lösas vid en definition av stadgan för grundläggande rättigheter .
Å andra sidan har vi också frågan om de sociala rättigheterna .
Här kommer det att bli nödvändigt att hitta en gemensam nämnare .
Å den portugisiska delegationens sida så skulle jag vilja säga att vi förstår att de ekonomiska och sociala rättigheterna är en del av Europeiska unionens arv som måste ingå i alla unionens dokument och i varje korpus med värderingar tillhörande Europeiska unionen .
Jag vet inte om den här uppfattningen delas av alla .
När det gäller den sista frågan så råder inte jämlikhet mellan män och kvinnor inom Europeiska unionen .
Jag är övertygad om att det här är en fråga som med största sannolikhet kommer att beaktas i stadgan , i synnerhet eftersom vi själva , när vi diskuterade Amsterdamfördraget , hade vissa uppfattningar om det , uppfattningar som sedermera fastslogs i Amsterdamfördraget varvid en kvalitativ förbättring gentemot Maastrichtfördraget uppnåddes .
Till sist och med anledning av stadgans införlivande i Fördraget om Europeiska unionen : Just nu leder jag den arbetsgrupp som vägleder regeringskonferensens beredningsgrupp .
Det är i portugisiska ordförandeskapets intresse att garantera att man efter ett godkännande av de personer som håller på att utforma stadgan - som ni vet så har rådet inte hand om stadgan , det ligger hos ett konvent med vald ordförande och med företrädare från Europaparlamentet , de nationella parlamenten , medlemsländernas regeringar samt Europeiska kommissionen - se till att det snarast blir färdigt ( det är fråga om ett förfarande som vi inte kontrollerar , som vi bara följer genom en vice ordförande från konventet som samtidigt är företrädare för Europeiska unionens ordförandeskap i samma grupp ) .
Det vore enligt vår mening önskvärt att stadgan införlivades i det nya fördraget för Europeiska unionen och att frågan genast remitterades till regeringskonferensen .
Jag tackar rådsordföranden för hans tankar och försäkringar om arbetets utveckling .
Ni förstår , min fråga har en mening , herr rådsordförande , eftersom rådet är ett av Europeiska unionens organ , och de europeiska medborgarna , såväl män som kvinnor , vill veta vilken dess vision är om Europas demokratiska och sociala modell i det 21 : a århundradet .
Jag skulle i min uppföljningsfråga vilja fråga er om ni , i egenskap av portugisiskt ordförandeskap , har planerat att barnens rättigheter - och här menar jag barnen som självständiga existenser - skall inbegripas i den diskussion som kommer att utvecklas och finnas med bland de rättigheter som kommer att införlivas i stadgan .
Fru talman !
Som sagt så har vi inte någon kontroll över själva utformningen av stadgan för de grundläggande rättigheterna .
Detta tillkommer de personer som ingår i den här gruppen och ärendet kommer bara att underställas rådet när och om man kommer överens om dokumentets lydelse .
När det gäller barnens rättigheter vill jag dock nämna att frågan är aktuell och har tagits upp av såväl Europeiska rådet som i en samling internationella dokument som vi har skrivit under .
Den här frågan skall tas med i stadgan för de grundläggande rättigheterna .
En fråga som min regeringen med all säkerhet kommer att driva inom ramen för stadgan för de grundläggande rättigheterna .
Vi har för övrigt även andra förslag .
Jag vet inte om förslagen i fråga kommer att godkännas eller inte .
Förmodligen är ämnet inte alltför polemiskt och det lutar åt en sammanställning av det som i dag är en samstämmig korpus för rättigheter som det inte vore mer än skäligt att inkludera i stadgan och delas av unionen .
Jag vill påminna ledamöterna om att frågorna , enligt anvisningarna till sammanträdet , skall vara koncisa och formulerade på ett sådant sätt att de kan besvaras i korta ordalag .
Ni känner till att parlamentet har en delegation med ledamot Méndez de Vigo som ordförande och ett utskott för konstitutionella frågor där dessa frågor kan diskuteras i detalj .
Därför ber jag att frågorna skall vara korta och likaså svaren .
I annat fall riskerar vi i viss mån att slå ut processen med framtagandet av en stadga om de grundläggande rättigheterna .
Jag ser att rådets tjänstgörande ordförande är villig att svara på allt , men min uppgift är att se till att frågestunden fortlöper .
Jag överlämnar ordet till Rübig .
Herr talman !
Fjorton medlemsstater har utlyst bilaterala sanktioner mot en medlemsstat därför att man där har bildat en demokratiskt vald regering .
Bägge partierna har redan suttit med i regeringen en gång .
Någon lagkränkning har det hittills inte varit fråga om .
Är förebyggande sanktioner förenliga med stadgan om de mänskliga rättigheterna ?
Vore det förenligt med stadgan om de allmänna fri- och rättigheterna om rådsordföranden gavs vetorätt för regeringsbildningen i medlemsstaterna ?
Är det förenligt med stadgan om de allmänna fri- och rättigheterna att uppmana till våldsdemonstrationer ?
Ärade kollega !
Som rådsordförande har jag inget svar att ge av den enkla anledningen att den ståndpunkt som intogs av den portugisiske premiärministern , som företrädare för fjorton statschefer och regeringar i medlemsländerna , gjordes bilateralt och inte i egenskap av ordförande i Europeiska unionen .
Jag vill dock påpeka att de förebyggande åtgärder som vidtogs på ett strikt bilateralt plan av Europeiska unionens medlemsländer har att göra med en rad åtgärder , som jag skulle vilja kalla profylaktisk politik på ett diplomatiskt plan , som vi menar är helt berättigade och rimliga när det gäller ett partis eller en partimedlems uppträdande i en regering i Europeiska unionen som inte verkar kunna garantera att unionens mål efterlevs .
Herr talman !
Jag har äran att vara ledamot i det konvent som utarbetar förslaget till stadga , så jag skall inte be ordförandeskapet spekulera över innehållet eller fråga huruvida det anser att konventet bör vara rådgivande eller huruvida det bör ha juridiska befogenheter .
Vad jag skulle vilja veta är vad som kommer att hända med det förslag till stadga som konventet utarbetar .
Kommer rådet att behandla det som ett dokument som det måste acceptera som det är , eller kommer rådet att känna sig fritt att ändra detta dokument ?
Kommer rådet helt enkelt att säga ja eller nej till det , eller kommer det i själva verket att ha möjlighet att sedan ändra förslaget till stadga ?
Svaret är varken ja eller nej .
Jag vet inte , ärade kollega , det beror på rådets beslut .
Fråga nr 8 från ( H-0042 / 00 ) : Angående : Beviljandet av exportkreditgarantier och de konsekvenser som detta får för byggandet av Ilisudammen i Turkiet .
Vid G8-mötet i Köln uppmanades OECD att inleda en process för att inrätta gemensamma standarder för beviljande av exportkrediter .
Dessa kan användas till att snedvrida konkurrensen och främja tvivelaktiga projekt .
Kommer EU att gå i bräschen för att denna process skall drivas framåt ?
Att det finns ett behov för detta framkom nyligen då den brittiska regeringen meddelade att den överväger att bevilja ett företag som deltar i bygget av Ilisudammen i Turkiet en exportkreditlicens .
Världsbanken har beslutat att inte finansiera projektet som kommer att innebära en omflyttning av 20 000 kurder , eventuellt en begränsning av Syriens och Iraks färskvattenförsörjning samt skador på miljön .
Vad anser rådet om det faktum att europeiska regeringar och företag deltar i detta projekt ?
Beträffande Caroline Lucas fråga så vill jag säga att man måste se på det ur två synvinklar : för det första exportkrediterna i allmänhet och för det andra vad som specifikt gäller för det här projektet .
När det gäller den mera allmänna aspekten så bör det påpekas att gruppen de åtta inte uppmanade OECD , som ledamoten insinuerar i sin fråga , att fastställa gemensamma kriterier för beviljandet av exportkrediter .
Kriterierna finns redan .
Avtalet som reglerar exportkrediter med officiellt stöd har varit i kraft inom OECD sedan 1978 .
Målsättningen med dessa direktiv är att se till att exportkrediter med officiellt stöd används på ett öppet och disciplinerat sätt .
De flesta OECD-länderna är som ni vet en del av det här avtalet , och Europeiska gemenskapen som sådan , inte medlemsländerna individuellt , är också en del av avtalet i enlighet med artikel 133 , före detta artikel 113 , i Fördraget om Europeiska unionen .
Avtalet har efterhand har ändratts och förbättrats , och Europeiska unionen vill fortsätta att vara gångjärn i den här processen eftersom det tycks ge oss större tyngd i de internationella ekonomiska förbindelserna .
När det gäller G 8 , och i enlighet med artikel 32 i uttalandet från toppmötet i Köln i juni 1999 , så har det sagts att vi tillsammans med OECD skall arbeta för att miljöfrågorna tas upp på ett likvärdigt sätt vid de exportbefrämjande institutionerna .
Vårt mål är att vara klara inför G 8-toppmötet år 2001 .
I G 8 är man alltså medveten om att det var det här som var det viktiga när det gäller exportkrediter och miljö och att det är det som OECD skall arbeta med .
I OECD : s ministerråd som jag deltog i 1999 välkomnade man de framsteg som hade gjorts när det gällde utarbetandet av ett OECD-avtal om miljöinformation för de större projekten vid exportkrediter med officiellt stöd .
Vi uppmanades också att fortsätta förstärka de gemensamma plattformarna under tiden som en rapport om de framsteg som gjorts färdigställs inför nästa ministerrådsmöte som äger rum i år .
Europeiska unionens medlemsländer har , som ni alla vet , en central roll i det här förfarandet och i den här diskussionen .
Mera konkret beträffande vattenkraftverket i Ilisu så förs samtal mellan de turkiska myndigheterna och de myndigheter vars exportkreditinstitutioner är potentiella leverantörer av kreditförsäkringar för export och projektets leverantörer som på ett tillfredsställande sätt bestämde sig för att värna om projektets miljömässiga , sociala och kulturella implikationer .
Det var för övrigt i det här sammanhanget som en företrädare från Förenade kungadömet i december 1999 tillkännagav att syftet var att garantera att exportkreditförsäkringarna underställs den typ av frågor som dem som ledamoten nämnde i sin fråga .
Frågan om exportkreditlicenser togs inte upp i samband med projektet .
Det bör påpekas att eftersom man inte har ansökt om lån för projektets finansiering av Världsbanken så riskerar man heller inget beslut om avslag från bankens sida .
Ett avslag kan man bara få om man har ansökt om något , förstås .
Det är tydligt att engagemanget från medlemsländernas regeringar och officiella exportkreditinstitutioner i vattenkraftverksprojektet i Ilisu fortskrider enligt de förpliktelser och det politiska och juridiska ansvar som länderna i Europeiska unionen , OECD och G 8 har tagit på sig .
Processen med att enas om dessa gemensamma standarder kan ha startat så långt tillbaka som 1978 , med det faktum att den brittiska regeringen tycks sätta igång med ett projekt som är väldigt skadligt för miljön antyder helt klart att den inte har varit särskilt framgångsrik hittills .
Jag undrar om ni skulle vilja svara på en fråga om investeringar av EU-företag i ansökarländerna .
Jag frågar detta med anledning av frågan om samstämmighet , ämnet för debatten i förmiddags .
Å ena sidan ber vi ansökarländerna att acceptera miljöregelverket , men ändå , på samma gång , stöder och uppmuntrar EU-medlemsstaterna investeringar i dessa länder som i sig själva är enormt skadliga för miljön .
Kan ni tala om huruvida frågan om investeringar i ansökarländer har förekommit i någon av de diskussioner fram till i dag som ni har hänvisat till eller inte ?
Ärade kollega !
Jag deltog inte i den debatt som ni hänvisar till .
Vad gäller den här delen av er fråga kan rådet bara besvara den skriftligt i efterhand .
Fråga nr 9 från ( H-0044 / 00 ) : Angående : Miljöproblem på grund av Drogheda Port Companys utvecklingsprojekt - revisionsrättens roll Det har uppstått en allvarlig konflikt mellan miljöskydd och strukturutveckling i området vid mynningen av floden Boyne i Irland .
Orsaken är ett utvecklingsprojekt som genomförs av Drogheda Port Company .
Det berörda området är ett särskilt skyddsområde enligt direktivet om vilda fåglar och man överväger för närvarande att klassificera det som ett särskilt bevarandeområde enligt habitatdirektivet på grund av dess internationella betydelse .
Många lokala och europeiska sammanslutningar har framfört hård kritik mot projektet .
Liknande fall förekommer i andra regioner i unionen : projekt som får EU : s utvecklingsstöd är inte ekologiskt hållbara .
Anser rådet inte att revisionsrätten bör ges ytterligare resurser i syfte att undersöka eller kontrollera dylika utvecklingsinsatser då det uppstår ekologiska konflikter ?
Vilka åtgärder ämnar rådet vidta för att stärka de europeiska institutionernas kontroll- och evalueringsbefogenheter i fall av denna typ ?
Med anledning av ledamotens fråga vill jag först och främst påpeka att revisionsrätten definieras i Fördraget om upprättandet av Europeiska gemenskapen .
I enlighet med artikel 246 i fördraget granskas räkenskaperna av revisionsrätten varvid alla gemenskapens inkomster och utgifter granskas , tillika regelbundenheten och legaliteten för nämnda operationer , dessutom står man som garant för en sund finansiell förvaltning .
För övrigt även i enlighet med artikel 248 .
Revisionsrätten förfogar därför från och med nu över alla instrument som behövs för att fullgöra sina skyldigheter .
Beträffande ledamotens förslag om att utöka revisionsrättens medel , anser rådet att alla unionens institutioner , inom ramen för gemenskapsbudgeten , förfogar över finansiella medel som gör att de på ett riktigt sätt kan verkställa sina respektive uppdrag .
I vissa fall hade det kanske varit önskvärt att utöka dessa medel men den möjligheten begränsas av budgeten , vilket ledamoten inte känner till .
Jag tar tillfället i akt och påminner om att Europeiska unionens budget gemensamt godkänns av rådet och parlamentet .
Rådet har därför inga möjligheter att ändra revisionsrättens uppdrag såsom det fastställts av fördraget .
Om extra resurser gavs till revisionsrätten , skulle det vara väl använda pengar , för det skulle säkerställa att EU-medel inte gavs till någonting som gick stick i stäv med våra miljöhänsyn .
Under flera år har rådet blockerat en bedömning av den strategiska utvecklingens konsekvenser hos projekt och program .
Jag skulle vilja fråga er om ni nu , när ni är ordförande i rådet , kommer att driva på detta ytterst viktiga förslag .
För det andra , eftersom det inte finns några hänvisningar till strukturfonderna i det nuvarande förslaget , skulle ni kunna se till de återinförs ?
Jag skulle vilja veta vad ni som rådets tjänstgörande ordförande kan göra åt detta just nu , för det är rådet som har blockerat detta under en lång tid .
Det är ytterst viktigt .
Om revisionsrätten regelbundet kunde bedöma de potentiella konflikterna mellan miljöhänsyn och strukturutveckling , skulle det vara mycket betydelsefullt , för revisionsrätten skulle kunna göra ett mycket värdefullt arbete .
Deras rapporter är utomordentligt detaljerade och mycket betydelsefulla .
Detta är ett sätt att se till att sådana konflikter undviks i framtiden .
Ärade kollega !
Många av era frågor faller under kommissionens behörighetsområde .
Det är följaktligen den som skall kontrollera vissa utvecklingsprojekts överensstämmelse med tillämplig miljölagstiftning .
Det är kommissionen som måste besvara de här frågorna .
Jag tror inte att jag kan ge ett bättre svar än detta .
Fråga nr 10 från ( H-0053 / 00 ) : Angående : Stadgan för Europaparlamentets ledamöter Rådet och Europaparlamentet skall försöka enas om en stadga för Europaparlamentets ledamöter .
En av de frågor som då skall regleras är om ledamöterna skall ha lika lön och var de skall betala sin skatt .
Enligt uppgifter i media anser det portugisiska ordförandeskapet att alla ledamöter skall betala samma skatt , till EU .
Detta står i strid med vissa medlemsländers uppfattning , vilka vill ha rätten att beskatta ledamöterna i hemlandet .
Kan det portugisiska ordförandeskapet klargöra sin position i frågan ?
Europeiska unionens portugisiska ordförandeskap är enligt min mening uppfylld av den här frågan .
Jag förmodar att det är första gången som man i ett arbetsprogram för ett ordförandeskap sätter upp och prioriterar problemet med Europaparlamentets ledamotsstadga på dagordningen .
Det portugisiska ordförandeskapet har därför sagt att man vill prioritera en lösning av stadgan , vilket för övrigt även Europaparlamentets ordförande sade vid Europeiska rådets möte i Helsingfors .
Vi är därmed i perfekt harmoni med varandra när det gäller att uppnå ett positivt resultat i den här frågan .
Det är med den här politiska viljan som vi försöker dra upp linjerna för en kompromiss och arbetet med detta har vi redan inlett .
Uppgörelsen måste nå enhällighet i rådet , vilket det är värt att påminna om , i enlighet med artikel 190 samt parlamentets bifall som måste godkänna stadgan .
Ordförandeskapet har inlett intensiva kontakter med flera av parlamentets ledamöter och med den grupp som parlamentet gav i uppdrag att förhandla med rådet .
Jag fick själv tillfälle att för första gången träffa gruppen under januarisessionen och jag tänker fortsätta med mina kontakter och träffa dem igen .
Debatten återupptogs av EU-rådets behöriga instanser , den här gången med större intensitet , och jag tror mig kunna säga att stadgans utformning är grundläggande för att samtidigt kunna garantera Europaparlamentsledamöternas självaktning och den nödvändiga öppenheten och sunda förvaltningen av allmänna medel , och detta säger jag i en anda där ökad flexibilitet råder och där vi alla är medvetna om hur viktigt det här är för allmänheten .
Beträffande den fråga som ledamoten ställde , vill jag påpeka att det inte är någon mening med en ny stadga om det inte innebär att situationen förbättras och ger dem som har identiska tjänster så likvärdiga villkor som möjligt .
Detta är utgångspunkten för det portugisiska ordförandeskapet .
Rollen som medlare tvingar oss dock att beakta alla åsikter som kan komma till uttryck i rådet och ledamoten är inte ovetande om att skattefrågan ställer till med problem i vissa delegationer .
I och med detta , och oavsett lösning , så menar jag att den demokratiska legaliteten alltid måste respekteras och accepteras av alla medlemsländer , oberoende av vad respektive nation har för åsikter .
Vad jag kan lova i den här frågan är att ordförandeskapet under sitt mandat kommer att arbeta i en anda av största möjliga genomblickbarhet och öppenhet gentemot ledamöterna och tillsammans med rådets ledamöter , i synnerhet dem som hade svårt att acceptera det förslag som dök upp förra året , så att man kan finna en rimlig kompromisslösning som samtidigt kan ge ledamotsstadgan den värdighet som behövs för det här huset .
Herr talman !
Jag tackar ministerrådet för svaret och vill ställa två följdfrågor som hänger samman med beskattningen av oss parlamentariker .
Min grundsyn är att man bör betala skatt i det land där man lever , där ens familj lever och där man har nytta av den offentliga servicen .
Jag tänkte fråga ordförandeskapet om det egentligen finns något argument för att vi inte skall betala skatt i våra hemländer precis som andra människor gör .
Finns det något argument för att vi skulle ha en speciell förmån därför att vi är just parlamentariker ?
Det är min första fråga .
Den andra frågan är om det portugisiska ordförandeskapet kan acceptera en lösning som innebär att skattefrågan löses på olika sätt för ledamöter av olika nationalitet , eller om ni vill ha en lösning som är lika för ledamöter av samtliga nationaliteter .
Ärade kollega !
Jag vill inte vara ohövlig mot kammaren , i synnerhet i respekt för ledamotens frågor , men låt mig slippa besvara frågorna punkt för punkt .
Vi är mitt inne i en ganska besvärlig förhandlingssituation , vilket visar sig i hur ordförandeskapet i Europeiska unionen ger uttryck åt något specifikt som har att göra med vissa situationer .
Detta drar givetvis med sig vissa konsekvenser då det bekämpas av andra ledamöter i rådet .
I den här fasen vill jag helst ursäkta mig och inte direkt besvara de frågor som ställs samtidigt som jag vill be er att döma oss efter de resultat som inom kort kommer att uppnås när vi försöker oss på en mera konkret lösning .
Jag kommer då gladeligen att inställa mig här i kammaren och besvara era frågor och förklara eventuella svårigheter om vi inte nått något resultat eller ta emot lyckönskningar av ledamöterna i fall resultat har uppnåtts .
Jag skulle vilja fråga rådets tjänstgörande ordförande om han , efter att under några få timmar här i kammaren ha arbetat tillsammans med dessa ledamöter av Europaparlamentet , har kunnat göra någon uppskattning av vad de är värda för lön ?
Ärade kollega !
Därför att den här debatten om Europaparlamentsledamöternas arvode inte bara är en debatt som berör ert land utan den berör även mitt land .
Jag vet exakt vilka arvoden som ledamöterna i Europaparlamentet betingar .
Jag är därför fullständigt medveten om problemet .
Herr talman !
Jag vill tacka för svaret .
Jag vill ställa en följdfråga som har en viss likhet med den Sjöstedt ställde .
Vi kommer båda från Sverige.I vårt land betalar vi vår huvudsakliga skatt i form av lokalskatt , eftersom servicen finns lokalt , och vi har en omfattande service .
Vi har problem med förtroendet för politiker , inte minst för europeiska politiker här i parlamentet .
Hur tror ni förtroendet för oss politiker skulle påverkas om det skulle bli så att vi får rätten att utnyttja servicen där vi bor - skola , omsorg osv - men samtidigt inte betalar någon skatt , inte bidrar ?
Hur tror ni ett sådant system skulle påverka förtroendet för oss politiker ?
Detta är en fråga , herr tjänstgörande rådsordförande , som jag inte är säker på att ni måste besvara , eftersom den är av filosofisk natur .
Men om ni vill ge er in på filosofiska resonemang , så varsågod !
Nej , herr talman , jag känner mig inte manad att gå in på filosofiska frågor .
Det här är frågor som berör grunden och har att göra med tanken bakom ledamotsstadgan och dess politiska roll .
Jag vill inte gå in i en sådan diskussion härför det verkar som om man då , för att använda ett franskt uttryck , à prejuger den tolkning som det portugisiska ordförandeskapet gör av förhandlingarna om ledamotsstadgan som man är inblandad i .
Eftersom tiden är ute för frågestunden med frågor till rådet kommer frågorna 11 till 35 att besvaras skriftligen .
Jag förklarar härmed frågestunden avslutad .
( Sammanträdet avslutades kl .
19.05 och återupptogs kl .
21.00 )
 
Tal av Tjeckiens president Vaclav Havel Herr president , mina damer och herrar ledamöter !
Å Europaparlamentets vägnar har jag den mycket stora äran att önska Vaclav Havel , Tjeckiska republikens president , varmt välkommen .
( Applåder ) Jag skulle också vilja hälsa fru Havel välkommen , som har tagit plats på åhörarläktaren .
Välkommen , fru Havel .
( Applåder ) Det är inte första gången vi välkomnar er här i parlamentet , herr president .
Ni har redan talat en gång i plenarkammaren i Strasbourg , för nästan sex år sedan , i mars 1994 , och många av oss har ett mycket starkt minne av det tillfället , de kolleger som var parlamentariker redan då .
Kort efter det att Maastrichtfördraget trädde i kraft uttalade ni er för en förstärkning av de europeiska värdena , för en europeisk etisk dimension och för att unionen skulle öppna sig för Central- och Östeuropa .
För många medborgare , och inte bara i ert land , personifierar ni därför detta värderingarnas Europa , för vilket vi ständigt uttrycker vårt engagemang .
Efter två val till Europaparlamentet och en ny viktig reform av Europeiska unionens fördrag , har unionens förbindelser med Tjeckiska republiken genomgått en ytterst dynamisk utveckling .
Ett associeringsavtal har trätt i kraft och en gemensam parlamentarikerkommitté EU-Tjeckien har inrättats .
1996 lämnade ert land in en officiell ansökan om medlemskap i unionen .
1998 inleddes slutligen de officiella medlemskapsförhandlingarna .
Den europeiska integrationsprocessen har , liksom utvidgningsprocessen , ökat i tempo på ett imponerande sätt sedan järnridåns fall .
Slutet för den konstgjorda uppdelningen av Europa inledde en ny epok .
I dag står vi inför en historisk utmaning och många framtidsutsikter för alla européer .
Herr president !
Ni är en viktig symbol för denna utveckling .
Ni grundade och undertecknade Charta 77 , en rörelse för försvaret av de mänskliga rättigheterna som företrädde och krävde grundläggande värden under en dyster period i ert folks historia .
För att ha försvarat människans frihet och värdighet dömde den kommunistiska regimen er till fem års fängelse .
Men ni förlorade aldrig hoppet och historien har gett er rätt .
Det är nu tio år sedan som " sammetsrevolutionen " krävde Havel i presidentpalatset .
Under tio års tid har ni som president först företrätt det demokratiska Tjeckoslovakien och sedan Tjeckiska republiken .
Försoningen med era grannar har för er varit , och är fortfarande , ett mål som ni har försvarat med stor kraft och uthållighet .
Ni är en första rangens europé .
I dag förbereder sig Tjeckien för att bli medlem av vår union .
Ni håller säkert med mig , herr president , och det har erfarenheten visat oss , att unionens utvidgningsprocess inte alltid är utan fallgropar , och det gäller för båda parterna .
Tjeckiska republiken måste göra stora ansträngningar för att uppfylla samtliga villkor för ett medlemskap .
Europeiska unionen måste å sin sida anpassa sina institutioner och politikområden inför utvidgningen .
EU har redan tagit ett stort steg framåt i samband med Agenda 2000 .
Följande etapp , dvs. den institutionella reformen , genomförs det här året i och med inledningen av den nya regeringskonferensen , där Europaparlamentet är en fullvärdig deltagare .
Vårt ansvar i egenskap av parlamentsledamöter är att se till att utvidgningsprocessen präglas av en maximal öppenhet och insyn , så att Europeiska unionens och Tjeckiska republikens medborgare en dag via sina valda företrädare skall kunna godkänna Tjeckiska republikens anslutning till Europeiska unionen .
Herr president !
Jag har det mycket stora nöjet att ge er ordet .
( Applåder ) Fru talman , mina damer och herrar ledamöter , mina damer och herrar !
Frågan om européerna besjälas av en europeisk identitet , vid sidan av ett medvetande om och en känsla av nationell tillhörighet , är en fråga som i dag ofta kommer upp på dagordningen .
Med andra ord : känner sig européerna verkligen europeiska , eller rör det sig snarare om en abstrakt idé , en teoretisk konstruktion som söker förhärliga en geografisk beståndsdel för att göra det till ett sinnestillstånd ?
Denna fråga väcks bland annat i debatten om vilken del av suveräniteten som nationalstaterna kan och bör överlämna till Europeiska unionens gemensamma organ .
Vissa menar att om den klart beprövade nationella tillhörigheten alltför snabbt trängs undan av en föga upplevd europeisk tillhörighet , ja som kanske till och med uppfattas som en chimär , kan det endast gå illa .
Så hur står det egentligen till med vår europeiska identitet ?
Om jag själv ställer mig den frågan på djupet ; hur europeisk jag känner mig och vad det är som förenar mig med Europa , blir jag först lätt överraskad : det är först nu jag ställer mig denna fråga , under trycket av vissa aktuella politiska frågor och förpliktelser .
Varför ställde jag mig inte den frågan för längesedan , under den tid då jag började orientera mig i världen och reflektera om den och mig själv ?
Betraktade jag min tillhörighet i Europa som ett rent yttre element , som inte var så viktigt , ett element som inte bör vara föremål för kval , eller till och med uppta mina tankar ?
Eller ansåg jag tvärtom att min europeiska identitet var något som kom av sig självt och inte förtjänar frågor , granskningar , följder ?
Den andra eventualiteten är mer trolig : allt som jag engagerat mig för har varit så naturligt europeiskt att det aldrig har fallit mig in att betrakta det som sådant .
Jag har helt enkelt inte sett poängen med att bedöma det på det sättet , och mer allmänt , att jag skulle förknippa mitt tänkande med någon kontinent .
Eller ännu bättre : jag har en känsla av att jag , när jag var ung , till och med skulle ha känt mig något löjlig om jag förklarade eller skrev att jag var europé , att jag uppfattade saker och tänkte på ett europeiskt sätt , eller till och med uttryckligen åberopade Europa .
För mig skulle det ha framstått som mycket patetiskt och förmätet ; jag skulle ha uppfattat det som en mer högmodig version av de nationella patrioternas patriotism , som alltid har besvärat mig .
Med andra ord : jag var så uppenbart och naturligt europeisk att jag inte ens reflekterade över det .
Och det gäller utan tvekan majoriteten européer : de är i grunden européer , men de inser det inte , betecknar sig inte som sådana och i opinionsundersökningarna förvånar de sig något över att behöva uttrycka sin europeiska identitet på ett tydligt sätt .
En genomtänkt europeisk samhörighet tycks inte ha en lång tradition i Europa .
Jag betraktar inte detta som något positivt och jag välkomnar med nöje det faktum att den europeiska identiteten i dag börjar anta en mer tydlig form i det stora havet med " självklara " begrepp .
Genom att ställa oss frågor om den , genom att reflektera och försöka definiera dess karaktär , ger vi ett viktigt bidrag till en förståelse för oss själva .
Detta kommer att bli avgörande i vår mångkulturella och multipolära värld , där förmågan att uppfatta vår identitet är ett första villkor för en god samlevnad med andra identiteter .
Om nu Europa hittills har ägnat sig ganska litet åt sin egen identitet , är det utan tvekan för att Europa med orätt har betraktat sig som hela världen eller åtminstone som något högre stående än resten av världen , och vi har därför inte känt ett behov av att definiera oss i förhållande till andra .
Med beklagliga konsekvenser , givetvis , för det faktiska beteendet .
Att bedriva ett reflektionsarbete om den europeiska identiteten innebär att man frågar sig vilken samling värderingar , ideal eller principer som begreppet Europa frammanar , ja vad det är som kännetecknar Europa .
Och mer än så .
Det betyder också att man bör göra en kritisk granskning av denna samling , vilket ligger i själva sakens natur .
Och således snabbt inse att många europeiska traditioner , värderingar eller principer kännetecknas av en stor tvetydighet och att de flesta av dem kan leda till helvetet om de överdrivs , utnyttjas eller missbrukas .
Om Europa nu träder in i självprövningens era betyder det att Europa har en önskan definiera sig i förhållande till andra , men också att man söker efter vad som är bra inom Europa , vad som är förlegat och vad som hör framtiden till .
När jag för sex år sedan hade den äran att för första gången tala i denna kammare , tog jag upp behovet av att betona den andliga dimensionen och betydelsen av den europeiska integrationens värderingar , och erkände min fruktan inför det faktum att det europeiska byggets andliga , historiska , politiska och civilisatoriska mening riskerade att döljas av tekniska , ekonomiska , finansiella och administrativa frågor , med risk för att allmänheten skulle bli helt förvirrad .
Vid den tidpunkten kunde mitt uttalande föra tankarna till en provokation , och jag var inte säker på om jag skulle bli utbuad i Europaparlamentet .
Inget sådant inträffade , men i dag kan jag med nöje konstatera att samma ord inte alls har samma provocerande karaktär .
Under de senaste tio åren har Europa genomgått en dramatisk utveckling - järnridåns fall , det ständigt mer uppenbara behovet av att utvidga Europeiska unionen , den allt snabbare ekonomiska integrationen och arsenalen av nya hot som har uppkommit med denna period - och alla dessa beståndsdelar har med nödvändighet fått Europeiska unionen att öppna sig för nya , mer intensiva självprövningar , för att definiera och på nytt söka efter de värderingar som håller den samman och ger dess existens en mening .
Man för ibland fram tanken att detta sökande kommer för sent , att den kulturella och politiska integrationen och självprövningen borde ha föregått den ekonomiska integrationen , med andra ord att man har börjat med slutet .
Jag tror inte att det är en rättvis bedömning .
Efter andra världskriget konfronterades det demokratiska Västeuropa med minnet av de två världskrigens fasor och faran för en expansion av det totalitära kommunistiska herraväldet .
Vid den tiden var det nästan onödigt att tala om värderingar att skydda .
De var uppenbara .
Det som krävdes var däremot att ena väst på ett så att säga tekniskt sätt , och det så fort som möjligt , för att förhindra att ny diktatur skulle uppkomma eller till och med breda ut sig , men också för att hindra gamla nationella konflikter från att blossa upp på nytt .
Detsamma gäller utan tvivel min europeiska identitet : eftersom den var så naturlig för mig under så många år , ja till och med årtionden , föresvävade det mig aldrig att åberopa den uttryckligen .
Allt som Västeuropa skulle skydda var så pass uppenbart , att man inte kände ett behov av att definiera , analysera , fördjupa eller omsätta det i olika politiska och institutionella realiteter .
Och på samma sätt som jag först nu frågar mig om jag känner mig europeisk och reflekterar över vad det betyder , har det senaste decenniets historiska händelser utan tvivel tvingat det under uppbyggnad demokratiska Europa att bedriva en fördjupad reflektion om själva grunden för dess enande och om sina mål .
De stora europeiska värderingarna - såsom de har formats av Europas andliga , politiska och stormiga historia och såsom andra delar av världen har anammat dem , åtminstone vissa av dem - är tydliga : respekten för den unika människan , hennes friheter , rättigheter och värdighet ; solidaritetsprincipen ; likhet inför lagen och rättsstaten ; skydd för alla etniska minoriteter ; demokratiska institutioner ; en uppdelning mellan den lagstiftande , verkställande och dömande makten ; politisk pluralism ; respekt för privat ägande och det fria företagandet ; marknadsekonomi och en utveckling av det civila samhället .
Den nuvarande formen på dessa värderingar speglar givetvis också ett stort antal europeiska erfarenheter under modern tid , som har gjort att vår kontinent har blivit en första rangens mångkulturella mötesplats .
Tillåt mig att uppehålla mig vid en av dessa grundläggande värderingar , av skäl som jag kommer att redogöra för .
Det handlar om det civila samhället .
I västvärlden , dvs. den euroamerikanska världen av i dag , utgör det civila samhället - ett öppet , decentraliserat och mångsidigt samhälle som är uppbyggt på tilltron till medborgarnas och deras många olika organisationers suveräna oberoende - den demokratiska statens bas och en garanti för dess politiska stabilitet .
När Europeiska unionen inom kort skall öppna upp sina portar för de nya demokratierna - vilket enligt min mening är ett centralt intresse för EU - är det mycket viktigt , om inte avgörande , att unionen hjälper till med att återuppbygga och utveckla det civila samhället i dessa länder .
Det var inte av en slump som den kommunistiska diktaturen , kort efter dess makttillträde , var så ivrig att med våld slita sönder det civila samhällets ömtåliga struktur för att slutligen omintetgöra det .
Det var för att de visste att de aldrig skulle få en verklig kontroll över folket så länge det civila samhällets olika strukturer , som byggts upp nerifrån , skulle fortsätta att fungera .
Det som blev kvar av det genuina civila samhället levde vidare och utvecklades i det direkta eller indirekta motståndet .
De europeiska värderingarna överlevde således i denna miljö , inte tack vare utan trots det politiska systemet .
Den spontana struktureringen av ett samhälle kan självklart inte föreskrivas ovanifrån .
Men man kan skapa en miljö och villkor som gynnar dess utveckling .
Stödet till de nya demokratierna bör därför ingå i ett större sammanhang , nämligen en varaktig fördjupning och förstärkning av det civila samhället i hela Europa .
Ju mer varierade , differentierade och sammanflätade de olika europeiska civila strukturerna är , desto större beredskap får de nya demokratierna för att ansluta sig till dessa , och desto fortare etableras principen om förtroende för medborgarna och subsidiaritetsprincipen , vilket möjliggör en förstärkt stabilitet i de här länderna .
Men det är inte allt : grundvalen för Europeiska unionen som överstatlig gemenskap kommer också att befästas .
Konkret sett medför detta , bland annat och framför allt , att vissa sociala solidaritetsplikter överförs till lokala myndigheter och icke-vinstdrivande organisationer eller offentliga organ .
Ju lägre den nivå är där resursfördelningen äger rum , desto öppnare och mer ekonomisk blir denna fördelning och desto bättre täcker den samhällets mest varierande behov - som är svåra att skilja från en central utgångspunkt - och desto mer genuin blir den sociala solidariteten , eftersom den blir mer tydligt förknippad med konkreta personer eller deras organisationer .
Medborgares , sociala gruppers , kommuners och regioners genuina solidaritet är således den bästa jordmånen för den solidaritet som endast kan beviljas av en enda enhet , dvs. staten .
Och i en så stor överstatlig enhet som Europeiska unionen , som måste fungera som ett solidaritetsinstrument , krävs det att dess medborgerliga grundval är än solidare , än rikare .
Europeiska unionens livskraft är därmed beroende av , bland annat och kanske främst , på vilket sätt medborgarna känner att de tillhör en europeisk medborgerlighet .
En växande medvetenhet om alla symptom eller uttryck för nationell egoism , främlingsfientlighet eller rasistisk intolerans borde naturligtvis utgöra en del av denna nya känsla av europeisk tillhörighet .
Den appeasement-politik som i München mynnade ut i en kapitulation inför det onda , är ett av den moderna europeiska historiens bittraste kapitel .
Denna erfarenhet manar till vaksamhet .
Det onda måste bekämpas när det ännu ligger i sin linda , och det räcker inte att det bara är regeringar som gör det .
Regeringarnas inställning borde vara ett resultat av medborgarnas attityd .
( Applåder ) Omsorgen om säkerhet är ett annat uttryck för den sociala solidariteten .
Detta är en uppgift för staten eller en överstatlig gruppering .
Europeiska unionen har påbörjat ett intensivt arbete med att utforma en ny säkerhetspolitik .
Denna politik borde utmärkas av förmågan att snabbt fatta beslut och lika snabbt omsätta dessa beslut i handling .
För mig är det en ytterst viktig faktor .
Det är för övrigt hög tid .
Den senaste erfarenheten i Jugoslavien säger oss mycket om den frågan .
Enligt min uppfattning var Natos intervention en relativt tydlig demonstration ur flera aspekter .
För det första kan , i förekommande fall , ett krav på att ingripa utanför Europeiska unionens gränser framtvingas av en respekt för livet , den mänskliga värdigheten såväl som omsorgen om den europeiska säkerheten .
Ju starkare mandatet bakom ett sådant ingripande är desto bättre , givetvis .
Men man kan tyvärr också föreställa sig en situation där det saknas ett FN-mandat , samtidigt som en intervention skulle gagna många människor , hela Europa och den mänskliga civilisationen i sin helhet .
Jag är inte säker på att Europa var beredd att ens helt nyligen konfronteras med så pass riskfyllda situationer .
Europa har utan tvekan en mycket större beredskap nu , åtminstone på ett psykologiskt plan .
Jag tror att Europa snabbt borde dra nytta av detta för att också göra materiella eller tekniska justeringar .
För det andra krävs det mycket större insatser för förebyggande säkerhetsarbete .
I Kosovo och i Serbien , liksom i Bosnien-Hercegovina och många andra områden i f.d.
Jugoslavien , hade tiotusentals människoliv och ett stort antal materiella tillgångar kunnat besparas om världssamfundet haft förmågan att reagera på ett lämpligt sätt tidigare , i konfliktens början .
( Applåder ) Trots alla vädjanden och alla varningar för eventuella eller hotande terrordåd hände tyvärr ingenting .
Möjliga och tänkbara skäl är bland annat omsorgen om de mest varierande särintressen och materiella intressen samt regeringarnas oförmåga att ta risker för den goda saken eller det allmänna intresset .
För det tredje spelade Förenta staterna i det här fallet den utslagsgivande rollen , och det är högst sannolikt att världssamfundet inte skulle ha vetat vad det skulle göra utan deras energi , och att vi än i dag hade fått bevittna den fasa som ledde fram till en intervention i Kosovo .
Men Europa kan inte förlita sig på Förenta staterna i all evighet , i synnerhet då det handlar om ett europeiskt problem .
Europa måste ha förmågan att besluta sig för en lösning och lösa situationen på egen hand .
I dagens värld , där små enheter på legitim väg sluter sig samman i form av internationella eller överstatliga gemenskaper , vore det otänkbart att Europeiska unionen fortfarande är en respektabel del av världsordningen men utan att kunna komma överens om ett sätt att försvara de mänskliga rättigheterna , inte bara på sitt eget territorium , utan också på det område där EU agerar , dvs. inom den sfär som en dag kan komma att tillhöra unionen .
Som jag sade för en stund sedan , anser jag att utvidgningen är ett centralt intresse för Europeiska unionen .
Tillåt mig att framhålla den övertygelsen , genom att peka på detta än en gång .
Det handlar kanske om erfarenheten hos en man som har genomgått 40 år av kommunistiskt förtryck , vilket föregicks av det nazistiska herraväldet , eller kanske om den särskilda erfarenheten hos en invånare i ett land beläget i Europas centrum , ett land som under seklens lopp har blivit en korsväg för olika andliga strömningar och europeiska geopolitiska intressen , kanske till och med den plats där mer än en europeisk sammandrabbning har sitt ursprung .
Detta har gjort mig bestämt övertygad om att Europa är den enda politiska enhet där säkerheten är odelbar .
Idén om två Europa som lever sida vid sida , idén om ett demokratiskt , stabilt och välmående Europa på väg att integreras vid sidan av ett mindre demokratiskt , mindre stabilt och mindre välmående Europa , är enligt min mening mycket bedräglig .
Den påminner om tanken om ett varaktigt sammanboende i ett rum , där ena halvan är översvämmad och den andra inte .
Hur mångskiftande Europa än må vara , så är det odelbart , och alla allvarliga händelser i Europa kommer att få konsekvenser och återverkningar på resten av dess territorium .
I egenskap av en unik politisk enhet , har Europa i dag en möjlighet som det aldrig har haft under hela sin stormiga historia : att organisera sig på ett i grunden rättrådigt och fredligt sätt enligt principen om jämlikhet och samarbete mellan alla .
Inga fler våldshandlingar som utövas av mäktiga gentemot mindre mäktiga .
I stället är det ömsesidig förståelse och allmänt samförstånd , hur besvärligt och hur lång tid det än tar att uppnå detta , som bör vara den främsta principen för såväl organisationen som stabiliteten i Europa under nästa årtusende .
Med Europa avser jag i det här sammanhanget kontinenten i sin helhet .
Vi vet alla att Europeiska unionens utvidgning bör åtföljas av fortsatta och djärva reformer av EU : s institutioner .
Jag är övertygad om att regeringskonferensen kommer att bidra med realistiska förslag som får Europeiska unionen att framskrida i rätt riktning .
Men jag tror inte att de institutionella förändringarna inom Europeiska unionen kan stanna vid detta .
Tvärtom ; enligt min uppfattning kommer det att bli starten för en mycket lång process , som kanske kommer att ta årtionden .
Denna process bör präglas av en ständig omsorg om att påskynda och förenkla beslutsfattandet inom Europeiska unionen och att göra det mer öppet för insyn .
Låt mig nämna två mer konkreta punkter som jag redan har tagit upp vid ett flertal tillfällen , och som i mina ögon skulle kunna bidra till att dessa mål förverkligas i en mer avlägsen framtid .
I första hand anser jag att Europeiska unionen förr eller senare bör förse sig med en koncis och tydlig grundlag som kan förstås av alla ...
( Applåder ) en grundlag som alla Europas barn kan lära sig i skolan utan problem .
Denna grundlag skulle innehålla två delar , som brukligt .
I den första skulle medborgarnas och de europeiska staternas rättigheter och skyldigheter formuleras , de grundläggande värden på vilka det enade Europa vilar samt det europeiska byggets innebörd och kallelse .
I den andra skulle Europeiska unionens viktigaste institutioner beskrivas , deras främsta befogenheter och ömsesidiga relationer .
En sådan grundläggande lag leder inte automatiskt till att den union som är sammansatt av stater skulle genomgå en radikal omvandling till en stor federal stat , en tanke som euroskeptikerna är besatta av , utan gör det bara möjligt för invånarna i det framväxande Europa att skapa sig en tydligare uppfattning om Europeiska unionens karaktär .
På så sätt skulle de bättre kunna förstå och identifiera sig med unionen .
( Applåder ) En av de viktiga frågorna , som ofta och med rätta tas upp i samband med unionens institutionella reformer , är frågan om vad man skall göra för att unionens små medlemsländer skall vara säkra på att de större länderna inte ser till att de hamnar i minoritet , samtidigt som man behöver ta hänsyn till de olika staternas storlek på ett riktigt sätt .
En möjlighet skulle kunna vara att upprätta en andra kammare i Europaparlamentet .
Den skulle givetvis inte väljas i direkta allmänna val , i stället skulle de olika parlamenten sända dit sina respektive företrädare , låt säga tre per stat .
Om den första kammaren , dvs .
Europaparlamentet av i dag , skulle återspegla de olika medlemsstaternas storlek , skulle den andra stärka jämlikheten mellan staterna : där skulle alla medlemsstater ha ett lika stort antal företrädare .
Mot den bakgrunden skulle exempelvis kommissionen inte behöva sättas samman enligt nationell tillhörighet , och de nationella parlamenten skulle bli involverade på ett mycket mer operativt plan .
Hur den institutionella eller den föreslagna reformen än utvecklas eller genomförs , finns det en sak som framstår som särskilt klar : en oenighet eller en avsaknad av samförstånd i institutionella frågor får inte bromsa utvidgningen av Europeiska unionen .
Skulle det bli så , finns det risk för att en alltför försenad utvidgning får oändligt mycket farligare konsekvenser än en eventuellt ofullbordad institutionell reform .
Mina damer och herrar !
Den tekniska civilisation som föddes på europeisk mark omfattar i dag hela vår planet och har blivit avsevärt påverkad av element ur den euroamerikanska civilisationen .
Europa har därför ett särskilt ansvar för tillståndet i denna civilisation .
Men detta ansvar får aldrig mer anta formen av en våldsam export av egna värderingar , idéer eller varor till resten av världen .
Nej , tvärtom , Europa skulle äntligen kunna börja med sig självt och tjäna som exempel , som andra kan men inte är tvingade att följa .
Hela den moderna uppfattningen om livet - som ständig tillväxt och materiella framsteg , grundat på den självsäkra människan som tar sig för universums herre - är den europeiska andliga traditionens dolda och beklagansvärda ansikte .
Denna uppfattning om livet förutbestämmer också den nuvarande civilisationens hotfulla karaktär .
Vem annars skulle kunna sätta upp ett starkt motstånd mot dessa hot , om inte vår del av världen , som satte igång rörelsen , ja kanske till och med vår civilisations fria fall ?
Vid denna brytpunkt i historien förefaller det vara Europas uppgift att bedriva ett djärvt reflektionsarbete om sitt tvetydiga bidrag till världen : att förstå att vi inte endast har lärt världen mänskliga rättigheter , utan att vi också har visat den Förintelsen ; att vi inte bara har fått världen att - andligt - förverkliga den industriella revolutionen och sedan den informationstekniska , utan också att vanställa naturen för att mångfaldiga materiella rikedomar , plundra den på dess resurser och förorena atmosfären .
Det gäller att förstå att vi visserligen har banat vägen för en oändlig vetenskaplig och teknisk utveckling , men att vi har gjort det till ett mycket högt pris : dvs. att vi har utmanövrerat en hel rad mycket viktiga och komplexa mänskliga erfarenheter som har formats under flera årtusenden .
Europa måste börja med sig självt .
Vi kan göra besparingar , införa fastetider och respektera - i enlighet med den bästa av våra andliga traditioner - den högre kosmiska ordningen som något som överskrider oss och respektera såväl den moraliska ordningen som dess konsekvenser .
Ödmjukhet , vänlighet , artighet , en respekt för det vi inte förstår , en djup känsla av solidaritet med andra , en respekt för alla olikheter , en vilja att göra uppoffringar eller goda handlingar som endast evigheten kompenserar - den evighet som observerar oss , i stillhet , tvärs igenom vårt samvete : dessa värderingar skulle kunna och borde vara det europeiska projektets program .
Europa har , helt eller delvis , det 20 : e seklets mest avskyvärda händelser på sitt samvete : de tvåvärldskrigen , fascismen och det kommunistiska totalitära systemet .
Under det senaste seklet har Europa också upplevt tre positiva händelser , även om alla inte bara kan tillskrivas Europa : slutet på det koloniala herraväldet över världen , järnridåns fall och början på det europeiska bygget .
Det fjärde stora uppdrag som väntar Europa är i mina ögon att försöka visa , genom sin blotta existens , att det är möjligt att avvärja den stora fara som vår motsägelsefulla civilisation utsätter världen för .
Jag skulle bli glad om det land jag kommer ifrån kunde delta i allt detta i egenskap av en fullvärdig partner .
( Kammaren gav stående talaren varma och långa applåder . )
Herr president !
Å Europaparlamentets vägnar vill jag verkligen tacka er mycket varmt för det starka budskap ni gav oss , kollegernas applåder vittnar om det .
Jag skulle vilja tacka er ; ni gör rätt i att påminna om att den nationella tillhörigheten är helt förenlig med en europeisk tillhörighet .
Och med utgångspunkt i er personliga erfarenhet visade ni oss att den europeiska tillhörigheten inte är något som kan förordnas , utan något som kommer spontant , naturligt .
Jag har antecknat era ord , och det är något som vi alla känner mycket djupt .
Vi kan konstatera att ni har förblivit trogen de principer som alltid har väglett er , som alltid har väglett era handlingar , detta engagemang för grundläggande värden .
Ni erinrade om det tal som ni höll 1994 och som ni själv beskrev som något provocerande , men det finns fruktbara utopier och vi har tillsammans kunnat titta tillbaka på den väg vi har tillryggalagt .
Och sedan skulle jag också vilja säga att ni på ett mycket bra sätt framhöll det civila samhällets roll och betydelse - inte endast i kandidatländerna , utan också i alla Europeiska unionens länder - för att återskapa medborgarnas förtroende , för att återge förtroendet för den sociala solidariteten , som vi behöver .
Och för att - kanske - sammanfatta det jag uppfattade som allra starkast i era uttalanden , det är att ni framför allt ville erinra oss om att det europeiska bygget vid sidan av dess ekonomiska aspekter var ett andens verk .
Vi har självklart en mycket stark önskan att fullfölja detta verk tillsammans med er .
Tack , herr president .
( Det högtidliga mötet avslutades kl .
12.40 . )
 
AVS-EU : s gemensamma församling Nästa punkt på föredragningslistan är årsrapporten ( A5-0032 / 2000 ) av Corrie för utskottet för utveckling och samarbete om resultaten av arbetet i AVS-EU : s gemensamma församling 1999 .
( PPE-DE ) , föredragande.- ( EN ) Herr talman !
Jag hade hoppats på att få presentera denna rapport klockan nio på morgonen i stället för klockan nio på kvällen .
Jag hoppas att antalet ledamöter i kammaren inte är en indikation på intresset för vårt utvecklingsarbete med utomeuropeiska länder .
Det är hur som helst det normala förfarandet att rapporten om AVS-EU : s församlings verksamhet presenteras för ledamöterna i detta parlament , och jag har den angenäma uppgiften att göra det i kväll .
Återigen kan jag rapportera att två mycket framgångsrika sammanträden har ägt rum , ett i Strasbourg och ett i Nassau .
På många sätt utgjorde detta slutet på en gammal era och början på en ny .
AVS-EU : s gemensamma församling är en unik organisation i världspolitiken .
Var annars möts 86 nationer för att diskutera frågor av ömsesidigt intresse ?
Sammanträdet i Strasbourg var det sista som leddes av Lord Plumb .
Med anledning av det enorma arbete som han har utfört under en svår period , utsåg den gemensamma församlingens presidium i Nassau honom till hedersordförande , och vi önskar honom all lycka efter hans pensionering .
De två sammanträdena har dominerats av förhandlingarna om en förnyelse av Lomékonventionen , och jag ser fram emot undertecknandet av en ny konvention och dess snabba ratificering av alla de berörda länderna .
Jag kommer ihåg att kommissionär Marin , vid den senaste delrevideringen då jag var föredragande , sade att den revideringen skulle bli den sista .
Men , han hade fel , och jag vill berömma Philip Lowe och hans lag , som har arbetat så framgångsrikt bakom scenen för att få till stånd en ny konvention under mycket besvärliga omständigheter .
Jag blev också mycket glad över att höra rapporten i förmiddags från kommissionär Nielson , som har arbetat outtröttligt för att utgången av förhandlingarna skulle bli den rätta .
Jag vill berömma honom särskilt för hans framgång .
Jag vill även berömma Kinnock och hennes arbetsgrupp för den enorma mängd arbete som de har lagt ned på Lomés framtid .
Jag är ganska säker på att Kinnocks rapport liksom rapporten om regionalt samarbete och integrering har haft stor betydelse för utgången av dessa förhandlingar .
Jag tackar även arbetsgrupperna för små östater och för klimatförändringar liksom gruppen för uppföljning av fisket för deras enastående rapporter .
Vi har haft frågestunder med rådet och kommissionen och med AVS-rådet , och jag skulle vilja tacka dessa institutioner för det intresse som de har visat för vårt arbete .
Det huvudsakliga målet med vårt arbete vid båda sammanträden gällde bekämpningen av fattigdomen .
I den antagna resolutionen gick man så långt som till att säga att fattigdom är liktydigt med en kränkning av de mänskliga rättigheterna .
I resolutionen betonades också betydelsen av att avskaffa ojämlikheter mellan könen , och när jag reser genom Afrika och ser det arbete som har utförts av kvinnor , önskar jag bara att det fanns fler kvinnor på högre regeringsposter och i presidentämbetet .
Vi skulle då kunna få se ett slut på en del av det bedrägeri , den korruption och den misshushållning som tycks vara endemisk i vissa länder och som måste stoppas .
Vi hade , som vanligt , många debatter om länder där det råder krigstillstånd .
Jag besökte Etiopien och Eritrea för att få förstahandsinformation .
Afrikanska enhetsorganisationen gör sitt bästa för att förhandla fram ett fredsavtal där .
Men Etiopien kräver fortfarande att vissa frågor skall klargöras , och den humanitära situationen i de båda länderna är allvarlig .
Vi blev i Nassau mycket glada över att höra att ett handelsavtal kan slutas med Sydafrika efter fyra års förhandlingar .
Detta belyser problemen med samstämmighet mellan EU och utvecklingsnationerna , något som fick sitt yttersta uttryck vid WTO-förhandlingarna i Seattle .
Det krävs mycket arbete för att övertyga utvecklingsnationerna om fördelarna med globalisering och världsomfattande frihandelsavtal .
I Nassau hade vi två intressanta debatter om Östtimor och Kuba .
Kuba har observatörsstatus , men jag förstår att landet nu har visat en vilja att ansluta sig till AVS .
Alla nationer som är belägna inom AVS-territoriets gränser och som kan leva upp till kraven på demokrati , mänskliga rättigheter , förvaltning av den offentliga verksamheten samt ett självständigt domstolsväsen är , är jag säker på , välkomna .
Jag avvaktar med intresse utvecklingen på Kuba .
När Dalmau , Kubas vice utrikesminister , talade inför församlingen , tvekade han inte att visa vilka känslor han hyste .
Angående Östtimor höll Da Costa , från Timors nationella motståndsråd , ett mycket rörande tal , i vilket han antydde att även Östtimor skulle vilja gå med i AVS när det blir en stat med en regering .
Vi måste ge dem allt vårt stöd för att nå det målet .
Mänskliga rättigheter är en så viktig fråga inom AVS-EU : s gemensamma församling att man har utnämnt gemensamma vice ordförande med särskilt ansvar för att på nära håll övervaka de mänskliga rättigheterna och rapportera till församlingen .
Ett antal fall har belysts , inklusive frågan om barnsoldater i Sudan , där många barn har blivit bortrövade från grannländerna .
Jag hade äran att bli vald till europeisk vice ordförande i inledningen av denna femte period , och Clair från Mauritius är AVS-ländernas nye vice ordförande .
Jag skulle vilja se ett antal förändringar i vår församling , särskilt efter undertecknandet av den nya konventionen i maj .
Vi måste få till stånd större jämlikhet mellan våra AVS-partner och våra europeiska medlemmar , och jag vill få ett slut på " de och vi " syndromet .
För det första skulle jag vilja se en gemensam parlamentarisk församling med valda ledamöter från AVS-länderna , i stället för att ambassadörer eller regeringsministrar sitter där som delegater .
Detta är , tror jag , den nya konventionen .
För det andra medges enligt den nya konventionen regionala församlingar i de sex regionerna , vilket skulle göra det möjligt för oss att vara mycket mer precisa i vårt arbete .
Dessa församlingar skulle rapportera till den gemensamma församlingen .
Vi hade en regional debatt i Nassau i Karibien , och den var utomordentligt produktiv .
Vi skall även hålla en debatt i Abuja i Västafrika .
Jag vill att församlingen skall upphöra med att vara enbart ett samtalsforum och i stället bli ett aktionsforum för förbättring av situationen för alla människor i utvecklingsländerna .
Jag vill att det civila samhället skall ges en högre röst .
Men för att det skall kunna göras , måste vi få ett slut på korruptionen , och vi måste angripa problemet rakt på sak .
Vi måste belöna de nationer som anstränger sig för att leva efter reglerna om god förvaltning av den offentliga verksamheten .
På samma gång bör vi slå ned hårt på dem som är korrupta eller vars författningar inte tillåter de pluralistiska regeringar som vi kräver .
Resultatet i Zimbabwe gör mig mycket glad .
De europeiska skattebetalarna kommer inte längre att acceptera att deras skattepengar används på ett otillbörligt sätt .
En ny vind av förändring måste blåsa över Afrika , och nya normer måste ställas upp och följas .
Den gemensamma församlingen bör spela en ledande roll när det gäller att övervaka tillämpningen av en god förvaltning av offentlig verksamhet , mänskliga rättigheter och demokrati i samarbete med kommissionen .
Jag tror att EU : s och AVS-ländernas valda delegater som likvärdiga partner klarar den uppgiften .
Jag ber att detta betänkande skall antas .
( Applåder ) Herr talman !
Låt mig först gratulera kollegan Corrie till det utmärkta och omfattande betänkandet .
Grunden för alla överläggningar om utvecklingspolitiken måste vara respekten för de mänskliga rättigheterna och kampen mot fattigdomen .
När fattigdom måste bekämpas så står minskningen av anslagen till utvecklingsbiståndet i många medlemsstater och i EU i skarp motsättning till detta .
Stickordet finansiering måste innebära att man med sikte på framtiden avsätter ytterligare medel för den gemensamma församlingen för att exempelvis kunna sända ut valobservatörer på begäran av AVS-länderna .
Vid samordningen av utvecklingsprojekten måste EU i framtiden för det första bli mer mångsidigt orienterad , för det andra komma bättre överens med de enskilda staterna för att arbeta effektivare och använda kapitalet på ett mer rationellt sätt .
Ett exempel vore utbildningen , som är det område där AVS-länderna i framtiden kommer att vara särskilt värda stöd och i störst behov av bistånd .
Om man då tänker på den rasande utvecklingen av möjligheter till utbildning och teknik via Internet så uppstår det helt nya hjälpmedel för att leda fram utvecklingsländerna med sina fortfarande blygsamma medel till globaliteten , inte globaliseringen .
Här ser jag en framtida uppgift för EU , nämligen att bidra till bildandet av en medelklass i AVS-länderna som är i stånd att fungera som hjälp till självhjälp .
Som exempel kan man titta på problematiken i Nigeria där man importerade färdiga produkter från industrin runt om i världen , men där underhållet kräver avsevärda kostnader för utländska hantverkare .
Lämplig utbildning av den nigerianska befolkningen skulle kunna bli vägledande för bildandet av en medelklass .
Den i rapporten tydligt utarbetade och absolut nödvändiga framtida optimeringen av arbetsmetoderna gör det , särskilt genom de tänkta regionala sammanträdena , möjligt att på ett bättre sätt ta sig an U-ländernas särskilda och olikartade problem , för vilka EU : s hjälpinsatser då kan förberedas mer målinriktat och sedan förverkligas .
Tack så mycket , herr Zimmerling .
Om jag är korrekt informerad så är det första gången som ni talar inför kammaren .
Det är ert jungfrutal , och jag skulle gärna vilja lyckönska er till detta .
Det gick alldeles utmärkt .
Herr talman , mina damer och herrar !
Det kan inte upprepas ofta nog : Loméavtalet utgör sedan 1975 en viktig stöttepelare för det europeiska utvecklingssamarbetet och innehar i många hänseenden en pilotfunktion .
I och med principen om partnerskap och paritet liksom att parlamentet har sällskap av den gemensamma församlingen är detta en världsmodell .
Lämpligt till jubileumsåret då vi får fira det 25-åriga Lomésamarbetet står vi inför att sluta ett nytt och mer utvecklat partnerskapsavtal som på bägge sidor också ger den gemensamma församlingen högre anseende som en äkta parlamentarisk församling .
Därför vill jag vid en tillbakablick inte inskränka mig till år 1999 ; det har föredraganden , Corrie , tagit ställning till på ett utomordentligt sätt .
Mycket av det som berör oss i dag är resultatet av grundläggande omvandlingsprocesser i alla delar av världen sedan slutet av 80-talet .
Detta har skakat om ordentligt även i U-länderna .
Efterskalven håller i sig .
AVS-samarbetet är en dynamisk process .
Från Lomé I till Lomé VI har det skett ständiga förbättringar av avtalsinnehållet .
Samtidigt har antalet partnerstater nu ökat väsentligt till 71 .
I synnerhet har utvidgningen kring Namibia och Sydafrika starkt berört alla som varit engagerade i frågan .
Nu har Kuba precis knackat på dörren , och om Kuba tas upp i AVS-EU : s gemensamma församling innebär det ett steg som får många konsekvenser och som inte heller låter sig tas utan förändringsprocesser på Kuba självt .
AVS-samarbetet förblir alltså högst spännande , inte bara på grund av de nya accentueringarna i det nya avtalet .
Fattigdomsbekämpning samt stödet till en hållbar ekonomisk , kulturell och social utveckling är viktiga målsättningar i arbetet med att i AVS-länderna bygga upp demokratiska samhällen som bygger på respekten av de mänskliga rättigheterna .
Detta inbegriper ett stärkande av de demokratiska institutionerna .
Här vittnar den gemensamma församlingens historia på ett imponerande sätt om en positiv utveckling .
Om det tidigare huvudsakligen var regeringsmedlemmar respektive regeringstjänstemän eller ambassadörer som satt kring bordet från AVS-ländernas sida så är våra samtalspartner i dag åtminstone till tre fjärdedelar valda företrädare från parlamenten .
Vi borde ställa till med en stor fest när det nu snart blir 100 procent , vilket ju är avsikten med det nya avtalet .
De fortskridande demokratiseringsprocesserna , som i motsats till de olika krisbildningarna i stor utsträckning löper obemärkt , uppmärksammas tyvärr alltför litet .
En specialitet i det multilaterala AVS-samarbetet är det regionala samarbetet respektive integrationen .
En önskning på Europaparlamentets långa önskelista kommer att uppfyllas : Den gemensamma församlingen kommer inom kort även att kunna hålla regionala sammanträden .
Detta har vi redan hört .
Ett starkare regionalt samarbete kan hjälpa till att förhindra att det bryter ut etniskt , ekonomiskt , socialt eller religiöst betingade konflikter , alltså ha en preventiv verkan .
Av samma anledning har Europaparlamentet sedan gammalt propagerat för att det civila samhället skall vara delaktigt i beslutsprocesserna liksom i ledningen för samarbetet samt framhävt betydelsen av ett decentraliserat samarbete .
De förstärkta kontakterna mellan den gemensamma församlingen och arbetsmarknadens parter som planeras i det nya avtalet är ytterligare ett steg i rätt riktning .
Återstår ett uns av motstånd i och med att den europeiska utvecklingsfonden fortfarande inte har lagts in i den europeiska budgeten .
Jag hoppas att det inte skall behöva ta ytterligare 25 år innan vi äntligen når resultat även här .
Herr talman !
Jag gratulerar herr Corrie till hans rapport .
Lomékonventionen har under 25 års tid varit ett uttryck för ett verkligt partnerskap mellan EU och AVS-länderna .
Att det överhuvudtaget har överlevt , trots det överväldigande motståndet mot det från många håll , inbegripet WTO , är en slags triumf .
Men den nya konventionen skall naturligtvis inte bedömas efter det faktum att den existerar , utan efter i vilken utsträckning den kan bidra till att EU : s åtagande att utrota fattigdom fullgörs och de internationella utvecklingsmålen nås .
Mätt med denna måttstock finns det ett antal allvarliga brister i de nya uppgörelserna .
Till exempel är avtalet särskilt misslyckat för de AVS-länder som lider av kortsiktiga svängningar i exportintäkterna .
Under ett maratonlångt förhandlingssammanträde i december nåddes en kompromiss , enligt vilken vad avser de minst utvecklade inlands- och östaterna , hjälp skulle ges i händelse av en minskning av exportintäkterna på minst två procent , i stället för vid den nivå på tio procent som gäller för andra AVS-länder .
Men vid det avslutande förhandlingssammanträdet hävdade EU att man i själva verket aldrig hade sagt ja till att inbegripa östaterna och inlandsstaterna staterna bland dem som skulle vara berättigade till stödet på grundval av tvåprocentströskeln .
Denna omsvängning har varit förödande för Winwardöarna i synnerhet , som kan vara det enda AVS-landet som faktiskt kommer att förlora kraftigt på de nya uppgörelserna .
Detta verkar vara en särskilt besynnerlig utgång , eftersom Winwardöarna är ett av de minsta och mest sårbara AVS-länderna , och de måste nu betala det högsta priset för denna nya Loméuppgörelse .
Under tiden , på handelssidan , har påtryckningar från WTO om att Lomékonventionen måste vara WTO-förenlig medfört att det finns en enorm kraft bakom idén med de så kallade regionala ekonomiska partnerskapsuppgörelserna eller frihandelsavtalen .
De länder som inte är bland de minst utvecklade länderna kommer med stor sannolikhet att utsättas för ett ansenligt tryck för att godkänna dessa uppgörelser .
Ändå är det ganska uppenbart att det även efter en övergångsperiod kommer att finnas ett antal länder som helt enkelt ännu inte kommer att kunna öppna sina marknader för frihandelns isvindar utan att den egna inhemska ekonomin ödeläggs .
Vi måste därför vara särskilt vaksamma och se till att det finns verkliga alternativ för de länder som inte ännu är redo för frihandelsuppgörelser .
Vi måste se till att strategier för att främja regional integrering inom AVS drivs efter egna linjer .
Avslutningsvis , under en eventuell ny handelsrunda bör EU och AVS-länderna gemensamt trycka på för en reform av GATT : s artikel 24 , för att uttryckligt erbjuda regionala icke-ömsesidiga handelsavtal mellan strukturellt och ekonomiskt olika grupper av länder .
Lomékonventionen är ett unikt partnerskap , men om det skall bli verkligt effektivt , måste det sträcka sig bortom diskussionerna inom Loméramen och inbegripa deltagande av WTO och ett partnerskap i alla andra internationella förhandlingsforum .
Herr talman !
I denna debatt vill jag kritisera den lott man tilldelar de fattiga länder i Afrika , Västindien och Stilla havsområdet som man vågar påstå är Lomékonventionens förmånstagare .
Inte ens på handelsområdet har Lomékonventionen på något sätt skyddat dessa länder ; deras andel i handeln med Europa har halverats , trots att den är obetydlig .
Detta återspeglar den ökade ojämlikheten mellan EU- och AVS-länderna .
Lomékonventionen tjänar framför allt några stora industriella eller finansiella företagsgrupper , som fortsätter att plundra dessa länder och upprätthålla deras ekonomiska beroende , särskilt i förhållande till de f.d. kolonialmakterna .
Det så kallade utvecklingsstödet tjänar uppenbarligen inte sitt syfte , eftersom underutvecklingen i de flesta av dessa länder fördjupas i stället för att dämpas , när det inte utgör en förtäckt subvention till europeiska exportindustrier .
Dessa stöd är i första hand manna för de befintliga regimerna , utan att befolkningarnas fattiga majoritet får några fördelar av det .
Och även om de delas ut på ett riktigt sätt , skulle de inte räcka till för att finansiera de mest nödvändiga infrastrukturerna på områden som hälsa , utbildning eller dricksvattenförsörjning .
Sedan flera år tillbaka minskar stormakterna dessa redan löjeväckande små stöd .
Höjden av cynism är när detta görs med förevändningen att de mänskliga rättigheterna inte respekteras eller att det finns korruption .
Men vem skyddar de regimer som främjar korruptionen , om inte de rika ländernas regeringar ?
Man blundar faktiskt för de som verkligen är korrupta , de stora oljebolagen , vattenleverantörerna och de offentliga företagen , som det trots allt skulle vara möjligt att gå hårt åt , eftersom de har sina huvudkontor här i Europa .
Debatten om valet mellan en förlängning av Lomékonventionen med dess kvoter och protektionism och en gradvis avveckling av Europeiska unionens och AVS-ländernas särskilda förbindelser i frihandelns namn , är en snedvriden debatt mellan två sätt att vidmakthålla plundringen och utarmningen av dessa länder .
Jag protesterar mot en simpel och omänsklig organisation som bokstavligen låter hundratals miljoner människor att dö i armod för att berika en minoritet .
Bara en obetydlig del av de enorma rikedomar som de stora företagsgrupperna har ackumulerat skulle göra det möjligt för dessa fattiga länder att ta sig ur misären , men så länge man inte vågar angripa dessa stora kapitalistiska grupper , döljer man bara problemen .
Herr talman !
Låt mig tacka ledamot Corrie , ordförande i AVS-EU : s gemensamma församling , som har haft den inte alltför avundsvärda uppgiften att sammanställa en rapport om en så svår församling som AVS-EU .
I detta mitt inlägg vill jag bara ta upp ett par punkter som jag anser vara av grundläggande betydelse .
Jag anser att Europaparlamentet med kraft måste kräva att församlingen verkligen blir parlamentarisk , dvs. uppmana AVS-länderna att låta sig företrädas av ledamöter från de nationella regeringarna , i syfte att förstärka AVS-ländernas demokratiska väv .
Låt mig i dag lämna mitt bidrag till debatten och peka på globaliseringen och den gemensamma organisationen av marknaden , som AVS-länderna ser som ett latent hot för den egna utvecklingen .
Jag anser det är nödvändigt med en övergångsperiod för AVS-länderna , men det är också nödvändigt att de får stöd mot bakgrund av de nya tankarna om en regionalisering av stödet , inte bara när det gäller jordbruket och fisket , utan också när det gäller utnyttjandet av gruvor och andra resurser under mark , av vilka några exploateras utan att AVS-länderna får annat än en blygsam ersättning .
Den tredje punkten gäller de ansträngningar som Europaparlamentet - via en gemensam arbetsgrupp inom ramen för den gemensamma församlingen - skall göra för att försöka stabilisera AVS-ländernas budgetar genom ett kvalificerat urval av budgetposter , för att möjliggöra en ekonomisk , men framför allt social , utveckling , och genom en övervakning av den inkomst- och skattepolitik som så småningom kommer att gälla inom AVS-länderna .
Vi måste stödja befolkningarna i AVS-länderna genom kontakter med deras regeringar , och de måste vara fullständigt på det klara med att utvecklingshjälpen från Europeiska unionen skall gå till folken och inte till de eventuella oligarkier som i vissa länder kontrollerar alla interna och externa resurser .
Den fjärde punkten , slutligen : förhindrandet av etniska konflikter och konflikter mellan olika länder måste vara en prioriterad fråga för oss och här kan man uppnå resultat såväl genom en kraftfull och auktoritativ diplomatisk offensiv som via de förslag som jag här har beskrivit .
Herr talman !
Jag ansluter mig till det positiva omdöme av rapporten som min kollega Karin Junker just har gett , och vill tillägga att Corrie har påbörjat sin uppgift som vice ordförande för den gemensamma församlingen AVS-EU genom ett effektivt och opartiskt agerande som verkligen förtjänar ett erkännande från vår sida .
Jag kommer att begränsa mitt inlägg till en viss händelse som ägde rum för bara några dagar sedan , delvis som en konsekvens av de händelser som tas upp i den rapport vi nu diskuterar .
Jag syftar på den önskan som Kuba gav uttryck för den 2 februari att som fullvärdig medlem ansluta sig till den grupp länder som bildar AVS .
En kubansk delegation deltog på AVS-EU : s senaste sammanträde i Nassau då vice förbundskansler Dalmau begärde ordet inför plenumet .
En livlig debatt utspelade sig som kom att följas av flera samtal mellan honom och många av oss .
Efter Nassau besökte en delegation från vårt parlament Habana under ledning av Corrie själv och Joaquín Miranda , ordförande för utskottet för utveckling och samarbete , och då ägde en rad klargörande åsiktsutbyten rum .
Jag har intrycket att delegationen från Europaparlamentet blev den sista påstötning som övertygade våra kubanska vänner om det lämpliga i att ta ett steg framåt mot ett samarbete med Europeiska unionen .
Vi befinner oss i en situation av stor politisk betydelse och jag hoppas att vi i Europaparlamentet kommer att skapa en ändamålsenlig och gynnsam vision samt visa en generös attityd från unionens sida i form av en snar positiv respons på Kubas ambitioner .
Det är viktigt , av minst tre olika anledningar .
I första hand för Kuba , för folkets utveckling och framgång och för att den blockad som införts av Förenta staterna en gång för alla skall hävas , en blockad som vid upprepade tillfällen har fördömts av Europaparlamentet och Förenta nationerna .
För det andra bör vi vara medvetna om att samtliga AVS-länder har uppmuntrat Kubas inträde .
Om vi från Europeiska unionens sida reagerar positivt på våra partners rekommendation , visar vi prov på respekt och hänsyn gentemot dem , något som kommer att vara positivt för vårt samarbete .
Man bör inte heller bortse från värdet av ett beslut som det jag föreslår , som bevis på Europeiska unionens samstämmighet och självstyre och på att vi inte är beroende av påtryckningar .
Genom att godta Kuba som medlem i AVS visar vi att Europa inte har fastnat i den hemska impulsen paying but not playing , och när vi protesterade mot vansinnigheter som lagen Helms-Burton gjorde vi det inte av skenhelighet utan för att vi är beredda att löpa linan ut .
Om några veckor kommer den gemensamma församlingen AVS-EU att samlas , och jag är övertygad om att den här frågan då kommer att behandlas .
Det vore önskvärt att Europaparlamentets företrädare i samband med detta stöder den kubanska strävan , så som parlamentskollegerna från AVS-länderna utan tvivel kommer att göra .
Kuba måste givetvis uppfylla de fastlagda villkoren på samma sätt som alla andra medlemmar .
Det vet kubanerna om och det åtar de sig garanterat att göra .
Det bör också klargöras att man inte kommer att begära mer av Kuba än det man har begärt av andra partner .
Vi välkomnar Kubas önskan om medlemskap och hälsar Kuba välkommet in i vår gemenskap .
Det säger jag helt uppriktigt men även utifrån en djup övertygelse om att , precis som blockaden inte har framkallat annat än elände och till följd av detta irritation och envishet från kubanernas sida , så kommer den integration som vi här stöder och den framgång som det leder till att ge upphov till det avspända läge och den öppenhet som vi alla vill ha och som vi alla , i synnerhet befolkningen på Kuba , kommer att ha nytta av .
Herr talman !
Jag vill också börja med att tacka och gratulera föredraganden , Corrie , för ett utmärkt betänkande som jag tycker väldigt väl beskriver och sammanfattar det arbete som har gjorts i AVS-EU : s gemensamma församling under 1999 .
Min talartid är kort , och jag vill egentligen bara ta upp två frågor : Den första frågan gäller fattigdomsbekämpningen som jag tycker börjar bli en pinsam historia både för EU och medlemsländerna .
Trots att man både i fördraget och på FN : s möten i Rio och Köpenhamn har förbundit sig att arbeta för att utrota fattigdomen i världen , skär man i själva verket ned på budgeten för utvecklingsstöd , tvärtemot vad man har sagt sig vilja göra .
Vi måste bryta denna trend .
Vi måste börja med skuldavskrivning .
Vi måste börja sätta aktion bakom orden .
Jag vill gärna att vi tar en ledande roll i detta arbete .
Den andra frågan gäller att vi i många sammanhang talar om att AVS-länderna måste lära sig demokratins grunder .
I punkterna 2 och 3 i resolutionen begär man inom ramen för den nya konventionen att arbetsmetoderna skall utvecklas och optimeras .
AVS-länderna skall uppmanas att låta många politiska opinioner komma till tals .
Det tycker jag är väldigt bra , och det skriver jag under helt på .
Vi måste emellertid också fråga oss hur vi själva hanterar demokratin .
Hur fungerar det inom Europaparlamentets delegation till AVS-EU : s gemensamma församling ?
I motsats till hur saker och ting fungerar här i Europaparlamentet och i parlamentets utskott , där man ju nominerar och utnämner föredraganden till betänkanden , finns det i denna delegation till den gemensamma församlingen inga som helst regler .
De två stora grupperna delar alla betänkanden , allmänna rapporter osv mellan sig .
För att ändra på denna odemokratiska ordning har vi , Verts / ALE-gruppen , lämnat in ändringsförslag 6 .
I detta ändringsförslag begär vi att föredraganden för betänkanden , och allmänna rapporter , samt medlemmarna i arbetsgrupper , skall utses enligt klara , demokratiska regler .
Hänsyn bör i detta sammanhang tas till små grupper och representativitet .
Herr talman , herr kommissionär , mina kära kolleger !
Jag vill i min tur först och främst gratulera vår kollega Corrie till hans utmärkta betänkande , som tydligt återspeglar debattinnehållet i den gemensamma församlingen , där han har varit en mycket effektiv vice ordförande .
Att utrota fattigdomen har stått i centrum för vårt arbete , och för att nå detta ambitiösa mål har många talare uppmärksammat kravet på att bevara ett mycket viktigt redskap , och då talar jag om förmånsavtalen mellan Europeiska unionen och AVS-länderna , inom ramen för Lomékonventionerna .
Detta är en stor utmaning .
Globaliseringen , avregleringen av handeln , WTO : s överhöghet och den internationalistiska filosofi som WTO förmedlar äventyrar själva kärnan i dialogen mellan Nord och Syd .
Man kan alltså bara glädjas åt att man har slutit ett nytt partnerskapsavtal för utveckling , och jag är för min del övertygad om att arbetet vid det senaste mötet i den gemensamma församlingen utövade ett avgörande inflytande för att få förhandlingarna att lossna , i likhet med det nya klimat som skapades efter händelserna i Seattle .
Jag gläder mig således åt att avtalen har förlängts , men det som framför allt fångar min uppmärksamhet är de nya vindar som nu blåser i våra förbindelser och som kommer till uttryck i den balanserade karaktären på de nyss avslutade förhandlingarna .
Europeiska unionen tycks äntligen ha brutit med den gamla paternalistiska logiken , och för att fatta mig kort , den neokolonialistiska logiken ; biståndsgivaren som gärna förvandlar sig till tillrättavisare , enligt en formulering som ligger vår vän Michel Rocard varmt om hjärtat .
Unionen har äntligen accepterat idén att ingen dialog är vare sig genuin eller effektiv om den inte antar formen av ett kontrakt som medför en respekt för respektive parts värdighet .
Genom att vägra lägga begreppet om god förvaltning i teknokraternas händer , så att det blir ett redskap för att skapa nya förbehåll , ger Europeiska unionen prov på klokhet och blygsamhet .
För oss tog det två sekel att lägga grunden till en demokrati vars skörhet vi ständigt blir påminda om i samband med aktuella händelser .
Med vilken rätt vill vi föreskriva vår modell för folk som ibland skiljer sig radikalt från oss i fråga om historia , värderingar och identitet ?
För min del föredrar jag den vilja som uttalas klart och tydligt i avtalen , dvs. önskan att öppna partnerskapet för nya aktörer - regionala myndigheter , icke-statliga organisationer - vilket för mig verkar vara den enda möjliga vägen för att successivt få dessa länders befolkningar att använda sig av samarbetet .
Att kort sagt gå från ett förödmjukande och infantiliserande stöd till ansvar , en garanti för effektivitet .
Herr talman , herr kommissionär , föredraganden , ärade kollegor !
Jag vill först och främst tacka för den exakthet och noggrannhet som ledamot Alexander Corrie har visat prov på i sin sammanfattning av betänkandet .
Europaparlamentets åsikt om AVS-EU-partnerskapet och dess aktiviteter , är oförnekligen av stor vikt för att nå politisk samstämmighet och befästa Europeiska unionens roll inom utvecklings- och samarbetsområdena .
Partnerskapets betydelse för bättre förbindelser mellan Europeiska unionen och AVS-länderna måste framhållas , ett partnerskap som blir alltmer parlamentariskt .
Inför en sådan positiv utveckling vore det i allas intresse att förse partnerskapet med en budget som är förenlig med ansträngningarna att göra ett kvalitativt arbete .
Inom ramen för partnerskapets verksamhet instämmer vi i föredragandens förslag att inrätta regionala parlamentariska församlingar i konventionens sex regioner , Karibien , Stilla havsområdet samt fyra afrikanska regioner .
Församlingarna skall följa aktiviteterna i respektive område .
Fattigdomen har varit den gemensamma nämnaren i alla partnerskapets debatter och utrotningen av denna det primära målet i Europeiska unionens utvecklingspolitik .
Kom ihåg att vi i enlighet med Nassaumötets resolution måste fullgöra våra åtaganden och minska fattigdomen såsom det internationella samfundet har beslutat .
Samstämmighet och handling är grundläggande .
Inför nästa Lomékonvention måste vi specificera hur mycket som skall investeras i utbildning , regionalt samarbete samt lokala myndigheters medverkan .
Det är mycket viktigt att lokal myndigheter kan medverka .
Samtalen om skuldsanering för de fattiga länderna genom program mot fattigdom och för en hållbar utveckling samt bekämpandet av bedrägeri och korruption är enligt min mening i ett vidare sammanhang grundläggande .
Vi måste gå vidare genom att vidta konkreta och samstämmiga åtgärder .
Befolkningen i de fattiga länderna börjar bli desperata .
Jag uppmanar kommissionen att vidta åtgärder för en snabb anslutning av Timor Lorosae till Lomékonventionen , så att man tillsammans med andra åtgärder kan bekämpa fattigdomen och påskynda den ekonomiska , kulturella och sociala utvecklingen och därmed förstärka den interna demokratin .
Avslutningsvis vill jag önska ordförandeskapet i rådet lycka till inför nästa toppmöte Europa-Afrika och be alla deltagare att arbeta för en konkretisering av de praktiska åtgärderna för befrämjandet av fred och demokrati samt utrotningen av fattigdomen i de afrikanska u-länderna . .
( DA ) Herr talman !
Jag vill gärna ta tillfället i akt och tacka föredraganden för det utmärkta betänkandet , och även tacka den gemensamma församlingen för dess arbete under 1999 .
Jag är också glad att kunna bekräfta att jag kommer att delta i den gemensamma församlingens nästa sammanträde som äger rum i mars i Nigeria .
Kommissionen vill att den gemensamma församlingen skall spela en större roll , särskilt när det gäller främjande av en bredare politisk dialog med våra utvecklingspartner .
Kommissionen håller med föredraganden om att kampen mot fattigdom även i fortsättningen skall vara det centrala målet för utvecklingspolitiken och att den alltid skall spela en nyckelroll .
Men för att det skall kunna ske en utveckling måste länderna delta aktivt i det globala ekonomiska systemet .
Vad gäller handeln med våra utvecklingspartner , är kommissionen helt inställd på att garantera att det vid varje nytt arrangemang tas hänsyn till AVS-staternas särskilda ekonomiska och sociala begränsningar .
Lucas nämnde att Stabex- och Sysminsystemet borde vara kvar .
Det håller jag inte med om .
Detta system har visat sig vara olämpligt , eftersom det faktiskt bara är till nytta för ett fåtal av de 71 länderna .
Det fungerar alltför långsamt och därför är det självklart att utvecklingsländerna accepterar det nya system som skall användas framöver , eftersom detta kommer att fungera mer flexibelt .
Jag kan med hänsyn till ländernas kommande anslutning till Lomékonventionen , som t.ex.
Östtimor , bara upprepa vad jag sade nyligen till Europaparlamentets utskott för utveckling och samarbete , dvs. att dörren är öppen .
Det är ansökarländerna själva som skall besluta om de vill knacka på dörren .
När detta skett tar vi ställning till det .
Kommissionen noterar vad gäller Kubas ansökan om tillträde till Lomékonventionen , att AVS-länderna enligt sin senaste förklaring stöder Kubas ansökan .
EU har alltid förespråkat en konstruktiv hållning gentemot Kuba , på samma sätt som uttrycks i EU : s gemensamma ståndpunkt , men det måste erkännas att diskussionerna kommer att bli komplicerade .
Rörande Elfenbenskusten kan jag informera om att alla 28 miljoner euro har betalats tillbaka i enlighet med vad som avtalats efter genomgången av de ekonomiska oegentligheterna .
Angående finansiering av Europeiska utvecklingsfonden över budgeten , kan jag säga att detta håller på att utvärderas .
Kommissionen stöder detta , men vi kan inte vid denna tidpunkt ge några nya rapporter om när eller hur .
Om artikel 366 a kan jag säga att det under förhandlingarna om ett nytt partnerskapsavtal fastställdes ett nytt förfarande för behandling av fall där det skett brott mot de mänskliga rättigheterna , de demokratiska principerna och rättsstatsprincipen .
Som det nu ligger till kommer parlamentet enligt Amsterdamfördraget på grundval av artikel 300 , att hållas fullständigt informerat om alla beslut och kommissionen kommer fortsatt att ta hänsyn till parlamentets resolutioner i denna fråga .
Det finns inga planer på att följa samtyckesförfarandet i parlamentet i samband med sådana beslut .
Det skulle nämligen kräva en ändring av det nyligen antagna Amsterdamfördraget .
Slutligen vill jag ta upp Sydafrikaavtalen , som föredraganden också tog upp .
Jag är helt enkelt glad - eller i det närmaste lycklig - för att jag här i kväll som en avslutning på denna debatt på ett mycket lämpligt sätt kan meddela att Sydafrikas president i dag har sagt ja till den lösning på de kvarvarande problem som rådet ( utrikesfrågor ) i måndags kom överens om att föreslå i samband med Sydafrika .
" Grappakrigen " är alltså slut .
Nu råder det fred och vi kan se fram emot ett samarbete med Sydafrika i enlighet med de gemensamma visioner och värden som denna fråga hela tiden egentligen skulle ha byggts på .
Jag tycker att det är en utmärkt grundsten för en debatt som i stort sett varit ganska positiv , och jag vill upprepa mitt tack till föredraganden och till parlamentet för det samarbete som sker med länderna i tredje världen i samband med just detta arbete .
Jag vill tacka er , herr kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Stabiliserings- och associeringsavtal med f.d. jugoslaviska republiken Makedonien Nästa punkt på föredragningslistan är betänkande ( A5-0031 / 2000 ) av Swoboda för utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik om rådets beslut om bemyndigande för kommissionen att förhandla om ett stabiliserings- och associeringsavtal med f.d. jugoslaviska republiken Makedonien ( SEK ( 1999 ) 1279 - C5-0166 / 1999 - 1999 / 2121 ( COS ) ) .
Herr talman , kommissionär Patten , kära kolleger !
Vi diskuterar i dag ett land som i sanning har genomgått svåra tider , ett land som dock med egna krafter , med egen vilja och säkert också med stöd av den internationella gemenskapen har utvecklats mycket positivt .
När Europeiska unionen , rådet och kommissionen , därför föreslår - och jag förmodar att parlamentet kommer att ansluta sig till förslaget i morgon - att det först och främst skall slutas ett stabiliserings- och associeringsavtal i Sydösteuropa , på Balkan - jag har inga skrupler att använda detta begrepp - då är detta i första hand ett tack eller ett erkännande för att på egen hand har arbetat sig fram till en bra position , ekonomiskt men förstås framför allt politiskt sett , med tanke på kriget i närheten och även i förhållande till den egna minoriteten .
Att utgöra en minoritet på 33 eller också 35 procent i det egna landet är med tanke på de omgivningar som landet befinner sig i nämligen inte någon bagatell .
Landet och dess politiker - säkerligen här och där i varierande grad - har alltid gjort ett gott arbete , och det skall erkännas .
Kommissionen föreslår att vi skall sluta ett avtal tillsammans med rådet .
Jag vill komma med ett par påpekanden , nämligen vad gäller just de områden där det måhända råder något differentierade uppfattningar , även om jag också här i särskilt hög grad vill lyfta fram och i berömmande ordalag nämna kommissionär Pattens arbete och intresse för och för hela regionen .
För det första : den regionala satsningen .
Jag anser att den regionala satsningen , om den förstås rätt , är både viktig och nödvändig .
Det måste finnas en beredskap för samarbete .
Så länge satsningen inte i viss mån uppfattas som tvång , utan som beredskap , som en möjlighet som borde utnyttjas av varje land , då är den riktig .
Det är bara det att när vi tittar på så ser vi att det i grannskapet finns en del länder som samarbetet t.ex. i ekonomiskt hänseende är mycket svårt med , som med Kosovo och Albanien , eller politiskt svårt som exempelvis med Jugoslavien .
Å andra sidan har samarbetet med Bulgarien och i synnerhet med Grekland utvecklats positivt , även det skall erkännas .
I detta sammanhang måste Europeiska unionen överväga - i början av veckan har man också börjat göra det - på vilket sätt grannlandet Jugoslavien - utan att man för den skull tar tillbaka något som helst av kritiken mot denna fruktansvärda regim - trots allt kan integreras i det regionala samarbetet .
Därför kommer jag i morgon att lägga fram ett ändringsförslag med vilket vi ställer oss bakom att sanktionerna koncentreras till regimen medan det å andra sidan ändå ges vissa lättnader för befolkningen och i den ekonomiska kooperationens anda även för näringslivet .
I detta hänseende - det får jag lov att säga eftersom jag kommer från ett land som Donau flyter igenom - är jag tacksam för de funderingar som kommissionen , dvs. kommissionär Patten har men även vice talman Palacio , som jag nyligen var i Budapest med , nämligen att göra Donau farbar igen för att möjliggöra ett minimum av ekonomisk återhämtning även för denna region , vilket självklart skulle vara mycket viktigt också för Rumänien .
Jag företräder uppfattningen att denna regionala satsning , om den förstås rätt , nämligen som ett sätt att bidra till den ekonomiska återhämtningen även på plats i själva regionen , är den rätta vägen .
Som sagt , som ett tvång får den inte uppfattas och heller inte ställas som villkor .
För det andra : Jag vill säga mycket klart och tydligt att vi vill att vägen in i Europeiska unionen skall stå öppen för och erbjudas .
Vi anser det vara en illusion att tro att det vore meningsfullt att yrka på medlemskap nu , men vi tycker också att det är fel att säga att det får vi tala om en annan gång .
Det är nu den vill ha svar på om man av princip kommer att ha denna möjlighet , när det väl är dags .
Landet fruktar att man så att säga skall utrangeras .
I hela omgestaltandet av stödverktygen ser man faran att inte längre vara sista vagnen på ett tåg som rullar i riktning mot Europa , utan att tåget skall köra vidare genom Europa medan man själv hamnar på ett uppställningsspår .
Men jag tror att kommissionär Patten har förståelse även för detta .
Jag ber honom eftertryckligen att klargöra också detta i lämpliga samtal .
För det tredje : Jag tycker att den - åtminstone hittills - också har visat sig vara i stånd att handskas bra med instrumenten .
Även om det naturligtvis krävs omställningar kommer den även fortsättningsvis att visa att många av de uppgifter som fortfarande i dag måste utföras i Bryssel framdeles kommer att kunna utvecklas i Skopje , i det egna landet .
Det är min förhoppning att mina kolleger skall kunna rösta för att vi godkänner dessa yrkanden som ett tecken på vår goda vilja gentemot den .
Herr talman !
Ända sedan krigen i Jugoslavien började har republiken Makedonien - jag använder helst detta förkortade namn - spelat en konstruktiv och fredsbevarande roll .
Vi erinrar om de förslag som regeringarna i Makedonien och då för tiden Bosnien-Hercegovina lade fram som syftade till att på ett fredligt sätt mildra och luckra upp den jugoslaviska federala strukturen .
Våra makedoniska vänner har således spelat en mycket positiv roll hela tiden , och av den anledningen måste det här sägas att Makedonien inte bara är ett objekt för vår så kallade stabiliseringssträvan , utan att det egentligen utgör ursprunget till denna .
Den förre presidenten Gligorov kan tillgodoräkna sig detta som en särskild förtjänst , och även den nuvarande presidenten har redan profilerat sig så mycket som president för alla makedoniska medborgare att Europeiska unionen inte kan göra annat än att skatta sig lycklig med en sådan samtalspartner på Balkan .
Trots alla anledningar som ligger för handen till eventuella nationella spänningar har de båda befolkningsgrupperna funnit en rimlig modus vivendi , och de fortsatta utsikterna till en ansvarsfull lösning av resterande problem är gynnsamma .
Tidigare var det framför allt i just Makedonien som jag hörde av romergruppen att de egentligen trivdes bra där .
Det hade jag inte hört särskilt mycket av romerna i Europa .
När det gäller problemen i Makedonien förtjänar den högre undervisningen för de albansktalande medborgarna särskild uppmärksamhet .
Tillgänglig högre undervisning , som man också har ett visst band till , är ett viktigt medel för att befolkningsgrupper skall kunna bli jämställda - det säger jag av egen erfarenhet som student vid ett protestantiskt universitet i Amsterdam .
Annars hade jag kanske aldrig studerat .
Ett sådant band och en sådan utbildning inom den högre undervisningen är också viktigt för utvecklingen av rättsstaten och även för de med rätta omnämnda lokala organisationerna , vilka måste förstärkas i sådana länder .
Avtalet med Makedonien måste också tillgodose en kompensation för den skada som landet ådrog sig på grund av den av oss beslutade bojkotten mot Serbien , som inte kostade oss något men Serbiens grannländer desto mer .
Om vi skulle kunna få en kursändring till stånd där skulle det vara positivt för oss med tanke på grannländerna .
Det är inte mer än rimligt att vi nu verkligen fastställer biståndet till Makedonien ordentligt .
Därför vill vi också ge vårt helhjärtade stöd till liberalernas ändringsförslag där man kräver att hjälpen inte skall bindas till givarländerna , för vi måste se till att biståndspengarna till återuppbyggnaden ger näringslivet i Makedonien och i regionen så många chanser som möjligt .
Där vill jag gärna räkna in Bulgarien och Rumänien också , för det förefaller mig vara ett taktiskt och psykologiskt fel att bara tala om de fem från före detta Jugoslavien plus Albanien .
För oss handlar det också om att ekonomierna i regionen kan stå på egna ben igen , vilket vi också har god möjlighet att få till stånd med biståndspengarna .
Avtalet med Makedonien måste kunna ses som att Europeiska unionen öppnar dörren för en anslutning av landet , även om detta fortfarande kommer att vara något på mycket lång sikt .
Under tiden måste vi i vår politik ständigt utgå ifrån hur önskvärt det är att Makedoniens lagstiftning verkligen börjar likna medlemsstaternas , och det måste återspeglas i vår politik , även i fråga om namnen på biståndsprogrammen för Makedonien .
Jag nämner här Phare-programmet som exempel .
Namnet på republiken , herr talman , är fortfarande ett problem på grund av att man är känslig för detta från grekiskt håll .
Jag utgår från att medlemsstaterna kommer att känna sig alltmer fria att på sitt eget språk använda den titel som passar för republiken .
Om vissa länder vill använda orden före detta Jugoslavien , då är det deras sak , andra behöver inte vara förpliktigade till detta .
Det handlar inte om att ständigt sätta oss under tryck .
Därför stöder jag Swobodas förståndiga betänkande ; vi hade inte heller väntat oss något annat av honom , och det är också anledningen till mina uppskattande ord om republiken Makedonien .
Herr talman , mina damer och herrar !
Låt mig först av allt personligen tacka föredraganden Swoboda för den utmärkta kvaliteten i hans arbete .
I dag uttalar vi oss positivt om att inleda förhandlingar om ett stabiliserings- och associeringsavtal med f.d. jugoslaviska republiken Makedonien .
Vi gör detta i medvetandet om att vårt beslut , det allra första som gäller detta område , innebär att en helt ny fas har inletts i våra förbindelser med Balkan .
Och avtalet är en del i denna nya fas , eller snarare denna politik som i en europeisk integration av regionen ser den enda möjligheten till en fredlig lösning av områdets konflikter .
Vårt bifall till förhandlingarna , så som dessa beskrivs i föredragandens motivation , uppkommer ur övertygelsen att det är rätt att i unionens politik kombinera såväl en regional dimension som ett mer specifikt utnyttjande av de ansträngningar som görs och de resultat som uppnås av de enskilda länderna vid anpassningen till gemenskapens acquis .
Det är denna dubbla målsättning som , enligt mitt förmenande , skall eftersträvas .
Å ena sidan skall man därför stödja de program som gäller till exempel infrastruktursatsningar , när man väl har förberett den tid - som ännu inte är inne - när vi kan se ett fritt handelsutbyte , efter att ha uppmuntrat de möjligheter som finns till ett ekonomiskt och kommersiellt samarbete mellan länderna i området och , å den andra , är det rätt att i dag tillsammans med f.d. jugoslaviska republiken Makedonien skapa förutsättningar för en politik som kan leda till en närmare integration .
För övrigt kan vår bedömning inte vara annat än positiv , av flera skäl .
Som vi har haft möjlighet att konstatera i våra besök till Skopje i den f.d. jugoslaviska republiken Makedonien , så har man gjort märkbara framsteg inom det ekonomiska området när det gäller demokratin och när det gäller en fråga som är mycket svår och omstridd på Balkan , den multietniska samlevnaden .
Å andra sidan är det pris man där har varit tvungen att betala på grund av kriget i det närbelägna Kosovo mycket högt , såväl när det gäller den praktiska hjälpen till Natos styrkor som när det gäller den minskade exporten till Nordeuropa .
Herr talman !
Låt mig avsluta med att bekräfta att dessa framsteg verkligen är vanskliga , bräckliga , osäkra och jag vill från vår sida uppmana till en konstant vaksamhet när det gäller de olika stegen i utvecklingen , steg som måste skiljas från varandra genom noggranna och regelbundna kontroller .
Herr talman , herr kommissionär , ärade kolleger !
Jag är här för att redovisa den värme och den hoppfullhet med vilken Europeiska liberala , demokratiska och reformistiska partiets grupp hälsar det faktum att förhandlingar inletts med den f.d. jugoslaviska republiken Makedonien .
Jag hyser gott hopp om att avtalet , inom de gränser som redovisats av föredraganden Swoboda , skall kunna bli ett föredöme , något som vi kan tillämpa i andra länder , framför allt Albanien , Bosnien-Herzegovina , Kroatien , Montenegro , Kosovo och , så snart som möjligt Serbien .
Vi är övertygade om att en snabb start för dessa förhandlingar och ett lyckligt slutförande av dem är den enda vägen om vi skall kunna nå fred i regionen - den fred som inte automatiskt följde när kriget i Kosovo tog slut - och att vi på så vis skall kunna undvika ytterligare sönderfall och att man återgår till kaos och våld , med alla de konsekvenser detta får vad gäller instabilitet för hela kontinenten , för att inte säga hela världen .
Om bevarandet av fred och säkerhet är det grundläggande motivet för den nuvarande djärva processen mot utvidgning av unionen till länderna i Östeuropa , så borde dessa motiv föreligga än tydligare i förbindelserna med Albanien och länderna i f.d. republiken Jugoslavien .
Detta kräver emellertid att man med beslutsamhet genomför den parallella utvidgning mot sydvästra Europa som nu sker genom de avtal som vi diskuterar .
Det är i denna anda , nästan som en provokation , som vi lagt fram ett ändringsförslag som skall överföra ansvaret för sydöstra Europa från utrikes frågor till utvidgningen .
Hoppet om att så snabbt och direkt som möjligt få med sydöstra Europa i de europeiska institutionernas arbete ligger bakom vårt förslag att även acceptera ett begränsat antal observatörer från de nationella parlamenten och Europaparlamentet och att personal från de aktuella länderna skall få arbeta inom domstolen och kommissionen .
För att uppmuntra regionens utveckling mot ett samhälle som är mer demokratiskt och bättre grundat på marknadsekonomiska principer är vi framför allt övertygade om att man måste göra omedelbara och konkreta framsteg för att intensifiera kampen mot korruptionen och göra den internationella hjälpen till återuppbyggnad och utveckling mer effektiv .
Därför har vi lagt fram ett antal ändringsförslag som vi hoppas att parlamentet skall acceptera : för det första att erbjuda den f.d. republiken Makedonien en tulltariff som motsvarar noll för exporten till Europeiska unionen och en kompensation för den progressiva minskningen av tullavgifter som Makedonien skall tillämpa på europeiska produkter , på villkor att man accepterar principen om en gemensam tullkontroll vid gränsen till Makedonien .
För det andra att den f.d. republiken Makedonien uppmuntras , genom lämpliga ekonomiska stödåtgärder , att gradvis koppla den egna valutan till euron som ett första steg mot en europeisering av hela den makedoniska ekonomin , dvs. med slutmålet att eliminera alla former av korruption från banksystemet .
För det tredje att den hjälp och det stöd som världen skall ge regionen , och därmed även Makedonien , skall vara tydligt multilateral till sin natur , utan att mottagarlandet får några direkta skyldigheter gentemot givarlandet .
Herr talman , ärade kolleger , herr kommissionär !
Vi hoppas att avtalet skall kunna uppfylla alla de mål som satts upp men vi skall inte inbilla oss att fred , stabilitet och välstånd i sydöstra Europa kan uppnås utan att man tar itu med betydligt större problem : jag tänker på Kosovos framtida konstitutionella status , nödvändigheten av att engagera Serbien i försoningsprocessen inom regionen och - varför inte ? - att åter diskutera förbindelserna mellan Europeiska unionen , Nato och FN , i ljuset av den nya balans som måste skapas mellan humanitära behov och statlig suveränitet , något som jag tror kommer att ändra strukturen för själva FN .
Herr talman , herr kommissionär !
Kosovokriget medförde att allting blev laddat .
Det gäller bestämt och framför allt för förbindelserna mellan Europeiska unionen och västra Balkan .
Sedan dess har förväntningarna varit högt uppskruvade .
Det gäller för situationen där , och det gäller för situationen här .
Där - eftersom man , vare sig vi tycker det är roligt eller inte , vid sidan av frågan om direkt stöd också ställer sig frågan : vad vill nu Europa med oss när allt kommer omkring ?
Finns det utsikter till medlemskap ?
Sådana frågor lever starkt i alla dessa länder .
Men även här är förväntningarna högt uppskruvade i Europeiska unionen .
Det första provet på om vi gör bra ifrån oss skulle kunna vara en äkta gemensam utrikes- och säkerhetspolitik .
Kan det lyckas för unionen att för första gången agera gemensamt och utveckla en gemensam politik för en så svår åtgärd ?
Det är också frågan om Europeiska unionen har lärt sig läxan av de dåliga erfarenheterna från Bosnien när det handlar om bistånd och de något bättre erfarenheterna från Kosovo .
Kan vi på grundval av erfarenheterna från Makedonien och fyra andra länder prestera ännu bättre ?
Mot denna bakgrund med mycket höga förväntningar tror jag inte att jag överdriver om jag säger att detta första steg , stabiliserings- och associeringsavtalet med Makedonien , är av avgörande betydelse .
Det är inte det enda bidraget från unionen .
Vi kommer inom kort till debatten om stabiliseringspakten , debatten om Cara-programmet och finansieringen på kort sikt .
Vi talar nu om stabiliserings- och associeringsavtalen , framtidsutsikterna på medellång sikt .
Därför tror jag att detta första avtal med Makedonien är så avgörande , för det är en förebild .
Jag är övertygad om att de andra fyra länderna kommer att fråga sig : vad kommer att hända ?
Vad kommer Europeiska unionen att göra med Makedonien ?
Kommer de att göra det som de gör med Makedonien med oss också ?
Det är på grund av att detta första steg fungerar som en förebild som det är så viktigt .
Makedonien är också en förebild i andra avseenden .
Föredraganden har redan påpekat detta på ett mycket klart och tydligt sätt .
Ta en sådan punkt som de interetniska relationerna .
Vi behöver inte återge detta på ett alltför idealiserat sätt här .
Vid presidentvalet visade det sig att det fortfarande inte står helt rätt till med allting , men jämfört med resten av regionen skulle man kunna tala om en makedonisk modell .
Det skulle vara mycket vunnet om vi tillsammans med makedonierna skulle lyckas att exportera den modellen till resten av västra Balkan .
Den förebildsmodellen gäller också för det regionala samarbetet .
Jag håller helt och hållet med föredraganden om att det där är nödvändigt att hitta en jämvikt mellan å enda sidan uppmuntran till regionalt samarbete och å andra sidan att bibehålla öppenheten till Bulgarien , till Grekland och att inte avskärma dem .
Herr talman , herr kommissionär !
Om vi lyckas bra med att ta detta första steg , då är väldigt mycket vunnet .
Om vi sjabblar bort detta , då är ännu mycket mer förlorat .
Herr talman !
Låt mig inleda med att konstatera att jag inte ser några problem med att principiellt stödja detta mycket väl underbyggda betänkande .
Jag vill bara peka på en fråga som enligt min mening saknas i betänkandet och som innebär ett stort problem för Makedonien och effektiviteten i ekonomiska och andra stöd från EU .
Jag talar om sanktionerna mot Jugoslavien .
För att undanröja missförstånd : Även jag anser att det behövs en effektfull uppgörelse med Milosevic-regimen .
Men för det första drabbar sanktionerna på ett omfattande och negativt sätt många av grannländerna , däribland Makedonien , som även utan detta befinner sig i en svår ekonomisk situation .
För det andra görs hela den jugoslaviska befolkningen genom underlåtenheten att respektera humanitära synpunkter på ett politiskt kontraproduktivt sätt ansvarig för Milosevic och hans krets .
Därför menar jag , vilket har formulerats i ändringsförslag 10 , att vårt ämne i dag borde föranleda oss att kräva ett snabbt slut på denna sanktionspolitik .
Herr talman , ärade kollegor !
Konflikten i Kosovo behövde inte avslutas innan vi kunde dra den slutsaten att det , efter flera krig i det forna Jugoslavien med de otaliga negativa konsekvenser detta förde med sig för stabiliteten i Balkan , är nödvändigt med en global och varaktig strategi för hela regionen så att fred och stabilitet kan garanteras i sydöstra Europa .
I den strategi som tog form genom den stabilitetspakt som antogs den 10 juni 1999 i Köln ser man regionen i sydöstra Europa som en helhet samtidigt som man också ser mångfalden och olikheterna i de länder som ingår .
Europeiska unionens bidrag till stabilitetspakten , till den så kallade " stabiliserings- och associeringsprocessen " , är ett exempel på utvecklingen av den regionala uppfattning som Europeiska gemenskapen utformade 1996 för regionens fem länder , Bosnien-Herzegovina , Kroatien , Förbundsrepubliken Jugoslavien , Makedonien och Albanien , vars viktigaste sida var fastställandet av politiska och ekonomiska villkor för att stödja fredsavtalet från Dayton , och därmed bidra till regionens stabilitet .
Att inleda förbindelserna mellan Europeiska unionen och Makedonien på en helt ny grund och öppna landet för en fullständig integrering i Europeiska unionens strukturer , genom det som förutsetts i stabiliserings- och associeringsprocessen , är av stor vikt för stabiliteten på Balkan .
Meningen är att länderna skall vara disponibla för ett godkännande av ett antal villkor .
Förhoppningen är att vi sänder dem en relevant politisk signal om att det en dag är möjligt för dem att bli en av oss , givetvis med respekt för deras egen suveränitet .
Efter att man erhållit vad som avtalats och utan några falska förhoppningar så kan det mandat som vi i dag är här för att ge kommissionen innebära det första stora steget mot fred och stabilitet i den så hårt plågade regionen , en region vars folk rättmätigt har visat att man vill tillhöra vårt område av frihet och utveckling .
Det är fullt tillräckligt med hur de fick lida under det sovjetiska oket och hur de sedan var tvungna att betala för att de hade tvångsintegrerats i det kommunistiska blocket .
Vi har informerats om att Makedonien ur politisk och ekonomisk synvinkel är berättigad att inleda nya avtalsförbindelser med Europeiska unionen , än mer efter det samarbetsavtal som trädde i kraft den 1 juni 1998 och som i praktiken reglerar respekten för gemenskapsarvet , i synnerhet på nyckelområden i den inre marknaden .
Mycket riktigt måste Makedonien fortsätta att uppbjuda alla sina krafter , men om man beaktar de politiska och ekonomiska reformer som redan har verkställts inom ramen för samarbetsavtalet och om man beaktar ett godkännande av övergångsperioder för vissa områden kan landet komma att uppfylla villkoren för ett avtal om stabilisering och associering .
Om vi utgår från tesen att landets utveckling är en stabilitetsfaktor för regionen , genom att definiera det föreslagna förhandlingsmandatet och genom att poängtera att det är fråga om ett bilateralt avtal med Europeiska unionen , så håller vi med föredraganden om att detta är den första konkreta tillämpningen av en långsiktig integrerad strategi för sydöstra Europa och att den fråga som ställs är att få veta hur Balkans strukturer på lång sikt skall se ut för att vara en garant för fred och stabilitet .
Ur ett sådant perspektiv blir syftet med ett regionalt samarbete grannländerna emellan i själva verket politiskt relevant .
Det här avtalet skall statuera ett exempel för de andra länderna i regionen .
Därför är det så viktigt .
Processen måste emellertid vara underställd en effektiv politisk vilja för ett närmande av de här länderna till Europeiska unionen .
Vi vet att ett av dem undergår en demokratisk stabiliseringsprocess , andra behöver fortfarande göra de demokratiska krafterna gällande i sina länder och andra uppvisar en jämvikt som är beroende av den militära närvaron i området , men det är länder som hädanefter vet att de , efter att ha överkommit svårigheterna , har en bro till sitt förfogande som kan leda till en effektiv förbindelse med Europeiska unionen .
Herr talman , herr kommissionär , kära kolleger !
Jag kommer inte att ansluta mig till mina kollegers kör av enhälliga röster .
Jag anser att detta betänkande är ett litet mästerverk i hyckleri .
I punkt 4 framhåller man hur föredömligt avtalet är .
Vi vet att det mellan Litauen och Turkiet finns 13 kandidatländer och att det finns en svart fläck i Europa , Balkan , och så vi vill få dem att tro att detta avtal är mirakulöst , samtidigt som vi förvägrar dessa länder möjligheten att vara kandidater .
I punkt 11 noteras att symboliska åtgärder kan ersätta det politiska avtalet , de politiska utsikter som erbjuds ett kandidatland .
Men det är inte bara ett mästerverk i hyckleri , det är också en absurditet , eftersom förhandlingarna påbörjas i morgon , kära kolleger , vilket innebär att avtalet kommer att undertecknas om ett år och träda i kraft om tre år .
Och då vill jag ställa er inför följande utmaning : finns det inte något land på Balkan som inom tre år kommer att lämna en ansökan om medlemskap i vederbörlig ordning - Kroatien , Makedonien , Bosnien ?
För några dagar sedan aviserade Racan att Kroatien kommer att lämna in en formell ansökan om medlemskap i slutet av år 2000 .
Jag är säker på att vi kommer att få fler ansökningar och då kommer detta fina arbete , denna vackra intellektuella arkitektur , att kollapsa , eftersom det kommer att bli förbisprunget av händelserna , precis om vi under 20 års tid har förbisprungits av allt som hänt i f.d.
Jugoslavien .
Detta skulle inte vara så allvarligt om det inte fanns de problem vi känner till i den här delen av Europa ; om det inte fanns de problem som man visserligen tar itu med , men som Makedoniens nya regering ännu inte har löst ; problemen med hur den makedoniska majoriteten och den albanska minoriteten skall kunna leva sida vid sida , med de nära sammanhängande problemen i Kosovo ; om det inte fanns de ekonomiska problem vi känner till , problemen med att bo granne med maffian , som är särskilt betydelsefull i Serbien ; om vi inte hade problemet med det veto som man absolut bör kritisera för vad det är , Greklands veto , som efter nästan tio år fortsätter att hindra detta land att kalla sig vid sitt eget namn , och jag hoppas att tolkarna inte använde termen FYROM ( före detta jugoslaviska republiken Makedonien ) när jag talade om Makedonien .
Detta är helt absurt .
Jag anser att det i första hand är en förolämpning gentemot våra grekiska kolleger , gentemot de grekiska medborgarna .
Den här frågan måste lösas så snart som möjligt .
Till sist har jag av en lycklig slump fått se ett brev som Georgievski , Makedoniens president , skickade till Fischler den 8 mars , där han frågar om Makedonien kan bli medlem av Europeiska unionen , med hänvisning till artikel O , i dag artikel 49 i fördraget .
Varför har inte rådet informerat oss ?
Varför har inte kommissionen informerat oss om denna formella begäran från Makedoniens sida ?
Herr talman , herr kommissionär !
Balkan är inte bara en mörk håla i politiskt hänseende .
Tänk på den påfallande positiva utvecklingen i Republiken Makedonien under de gångna , kritiska åren .
Den fruktansvärda etniska upptrappningen i det närbelägna Kosovo spreds inte till makedoniskt territorium .
Paradoxalt nog , men likväl sant , hade kriget på Trastfältet , Kosovo Polje , rakt motsatt effekt : en påtaglig minskning av den farofyllda förtroendeklyftan mellan den makedoniska befolkningsmajoriteten och den albanska minoriteten .
Ur de förstnämndas synvinkel uppförde sig de senare lojalt gentemot den gemensamma staten när Kosovokonflikten exploderade internationellt .
Och enligt den albanska minoritetens synsätt uppfyllde makedonierna liksom den makedoniska staten på ett frikostigt sätt sina förpliktelser gentemot den ytterst plågade albanska befolkningsmajoriteten i Kosovo .
Denna anmärkningsvärda konsekvens av krigshandlingarna i Kosovo kan därför med rätta kallas det andra , inre statsgrundandet av Republiken Makedonien .
Swobodas balanserade , aktningsvärda betänkande ansluter på ett mycket konkret sätt till detta överraskande och samtidigt glädjande resultat .
Kort sagt , Europeiska unionen vet vad den har att göra i Makedonien .
Hjälp denna färska tillflyktsort för mängder av krigsflyktingar att på ett tillbörligt sätt uppfylla sin roll som drivkraft för den tilltänkta stabilitetspakten på Balkan .
Herr talman !
Sedan åtta år tillbaka befattar jag mig med Makedonien , och jag vill gärna säga emot Dupuis .
Det är inte hyckleri vi ägnar oss åt .
Vi har kommit fram till en gynnsam tidpunkt , och jag tror att makedonierna uppskattar det .
Var nu inte stygg och häll vatten i deras vin .
Jag tycker att vi bör närma oss detta på ett mer positivt sätt .
Makedonien har inte varit i krig .
Men landet har lidit av kriget i omgivningarna och av sanktionerna , och det lider fortfarande av de sanktioner som med rätta har vidtagits mot grannländerna .
Man har lidit oändligt av flyktingströmmarna under Kosovokriget .
Därför måste man också säga att utvecklingen i Makedonien har löpt förvånansvärt kontinuerligt demokratiskt .
Det är ett land som inom sig har svåra interetniska problem att få bukt med och som också löser dessa på ett alltmer framgångsrikt sätt .
Jag vill tydligt poängtera att vi kan lyckönska Makedonien till en förebildlig minoritetslagstiftning och tillämpningen av denna , samt att det konsekventa inbegripandet av den 30 procent stora albanska befolkningen i regeringens agerande , i regeringspolitiken och i samhället är en förutsättning för den fredliga samexistensen i Makedonien .
Det gläder mig att den önskan som Swoboda har framfört i sitt betänkande kommer att gå i uppfyllelse i början av mars , dvs. att EU-delegationen där nere äntligen bildas , att vårt anseende som Europeiska unionen äntligen höjs där nere .
För mig är starten på förhandlingarna om stabiliserings- och associeringsprocessen den logiska slutledningen av en produktiv och god utveckling i landet .
Inom ramen för vårt politiska engagemang måste Makedonien äntligen få erfara i praktiken att dess eget glädjande regionala samarbete belönas även av oss genom att vi faktiskt drar igång regionala projekt .
Jag skall endast nämna två små : Den snabba lösningen på problemet vid gränsövergången till Kosovo i Blace och förverkligandet av korridor 8 , dvs. från Albanien via Makedonien till Bulgarien .
Jag anser att Swobodas betänkande är utomordentligt bra , och jag instämmer helt och fullt .
( Applåder ) Herr talman !
Jag skulle även från min sida gärna vilja framföra komplimanger till kollega Swoboda för hans betänkande .
Jag tror att det är bra att vi är så många här som uttalar stöd för den taktik som han väljer där .
Det handlar om att ta itu med stabiliteten i regionen på ett strukturellt sätt , och det är också innebörden i det kommande avtalet med republiken Makedonien som vi behandlar i dag .
Medan stabilitetspakten fortfarande väntar på det faktiska genomförandet har kommissionen mycket snabbt arbetat med att utveckla det nya instrument som heter stabiliserings- och associeringsavtal .
Därmed påbörjas arbetet med att fördragsmässigt stabilisera länderna i före detta Jugoslavien .
Det handlar om länder som ännu inte kan komma i fråga för ett föranslutningsavtal .
Det avtal som ligger framför oss är egentligen ett slags " före-före " , men då med möjlighet till framtida medlemskap .
Att på detta sätt binda länder via aktiva fördrag är ett utmärkt instrument under förutsättning att de avtal som fastställs där tillämpas fortlöpande för att den önskade stabiliseringen också skall uppträda .
Makedonien är fortfarande en potentiell krutdurk och har en historia som sådan .
Landet har dock ambitionen att bli befriad från denna beskrivning .
För detta syfte behövs inre stabilitet .
Den nya regeringen vill vara öppen för detta , och avtalet kan fungera som en dagordning för reformer , inklusive en direkt roll och en likaberättigad ställning för den albanska minoriteten .
Landet behöver nu framför allt lugn för att bringa ordning internt och finna vägen mot en större välfärd .
Vi , i synnerhet socialdemokraterna , vädjar till oppositionen att iaktta dessa uppfattningar .
De måste vara med och stödja den makedoniska modell som här lovordats så mycket .
Men landet behöver också och framför allt yttre stabilitet .
Vad tjänar inre stabilitet till om omgivningen är instabil ?
Denna stabilitet är nödvändig i förbindelserna med Jugoslavien , Kosovo , Albanien och Bulgarien .
Regionen måste erkänna att Makedonien existerar , och det kommer landet att fortsätta göra .
Yttre stabilitet innebär öppna gränser och regionalt samarbete .
Minoriteter och majoriteter måste få utrymme för mänskligt och kulturellt utbyte .
Stabiliteten i Makedonien hänger starkt samman med utvecklingen i grannländerna .
Kosovoproblemet är känt ; där finns världssamfundet närvarande i stor omfattning .
Det förefaller som om faktorn Albanien underskattas .
Unionen anser att tiden ännu inte är mogen för ett stabiliserings- och associeringsavtal med det landet .
Men vad skall det då bli ?
Det är just argumenten för att sluta ett avtal med Makedonien och att ännu inte göra det med Albanien som skapar så stark oro hos oss att en avvaktande hållning från unionens sida beträffande Albanien egentligen inte är godtagbar .
Hur hanterar kommissionen denna avvägning ?
Jugoslavien är i lika hög grad en svag stabilitetslänk och därigenom ett hot mot ett stabilt Makedonien .
Vi måste avvakta vad som sker där .
Stämningen i Belgrad blir allt mer oförutsägbar för varje dag .
Vi stöder emellertid rådets beslut att ge sanktionerna en annan betoning .
Det innebär i alla fall att vi äntligen gör ett seriöst försök att ge oppositionen , som förbereder sig inför en ny omgång demonstrationer , stöd i ryggen .
Vad skall unionen göra mer i den riktningen för att oppositionens krav - tidigarelagda val - skall infrias ?
Vad mer kan vi göra och företa oss för att stödja denna opposition ?
Herr talman , herr kommissionär !
Kosovo blev förhoppningsvis det sista fallet då folkrätt kunde tolkas som att diktatoriska ledare kunde förfölja minoriteter på det mest vidriga sätt med hänvisning att " det sker inom den egna nationen " .
När USA och Nato samt till slut också EU reagerade var det sent , mycket sent .
Mycket lidande hade kunnat undvikas om bl.a.
EU hade agerat tydligare och tidigare .
Vi , Europeiska unionen , har därför ett särskilt ansvar för att nu hjälpa , bistå och bygga upp Balkan .
Vår absoluta målsättning måste vara att skapa förutsättningar för alla länder i Sydösteuropa att integreras med övriga i EU - ekonomiskt , handelsmässigt och politiskt .
Att ge grogrund för demokrati i denna krigshärjade del av Europa sker bäst genom handel och ekonomisk integration .
Vi liberaler är beredda att gå långt och göra det fort , precis som Paolo Costa har redovisat .
Vi hälsar därför med största tillfredsställelse det förslag till stabiliserings- och associeringsavtal med Makedonien som nu föreslås och tackar Swoboda för ett mycket bra betänkande .
Makedonien förtjänar vårt stöd , inte minst med tanke på det uppoffrande , oegennyttiga arbete som Makedoniens befolkning och dess ledare visade upp under Kosovokriget .
När Makedonien nu sliter sig ur kommunismens och nationalismens förödande garn , är det vår skyldighet att mycket tydligt agera och stödja .
Precis så skall vi göra för de övriga länderna på Balkan .
Det är en bjudande plikt för EU .
Herr talman , låt mig i detta sammanhang påminna ledamöterna - inte minst med tanke på en diskussion tidigare i kväll - om att den man som bär huvudansvaret för krig , mänsklig förnedring , mördande och fördrivning av oskyldiga människor från deras hem fortfarande styr rest-Jugoslavien , Serbien .
Den man som är anklagad för folkmord och borde ställas inför krigsterminalen i Haag går fortfarande fri .
Jag talar om Milosevic .
Så länge som Milosevic är kvar och Serbien inte går en demokratisk väg , så länge utgör Serbien ett ständigt hot för freden på hela Balkan - också för Makedonien .
Herr talman !
Detta avtal kommer att utgöra den första tillämpningen av stabilitetspakten i sydöstra Europa .
Helt klart är att avtalets villkor , som godtas i Swobodas betänkande , inte har freden som mål , utan en större politisk och ekonomisk styrning av landet , kontroll över dess naturtillgångar , hård exploatering av dess arbetskraft och ytterligare utnyttjande av landet som bas för operationer mot de länder och folk i regionen som motsätter sig den nya ordningen .
Och allt detta i utbyte mot ett löfte om en framtida anslutning till Europeiska unionen .
I betänkandet godtas dessa riktlinjer , liksom Europeiska unionens allmänna politik för sydöstra Europa .
Det är betecknande att man i betänkandet ger komplimanger till före detta jugoslaviska republiken Makedonien ( FYROM ) för den konstruktiva hållning som landet intog under Natos attacker , man lovordar landets fredsfrämjande roll , eftersom det accepterade att Natostyrkor utplacerades på dess territorium ; naturligtvis tystar man ned folkets vrede , som kom till uttryck i omfattande protestaktioner under Natos bombningar .
Avslutningsvis , eftersom vi anser att såväl stabilitetspakten som det stabiliserings- och associeringsförfarande som Europeiska unionen tillämpar för länderna i regionen kommer att skapa nya problem i regionen , nya vedermödor för folken , liksom de kommer att stärka de amerikanska och europeiska imperialisternas dominerande roll ytterligare , kommer vi att rösta emot betänkandet och på så sätt ge uttryck för vår solidaritet med folket i den före detta jugoslaviska republiken Makedonien .
Herr talman !
Herr kommissionär !
Ett av de mest grundläggande målen för stabiliserings- och associeringsavtalet mellan Europeiska unionen och före detta jugoslaviska republiken Makedonien ( FYROM ) är att befästa stabiliteten och freden i regionen , något som naturligtvis förutsätter att goda grannförbindelser mellan de berörda länderna utvecklas och bibehålls .
Jag skall inte uppehålla er med detaljerna i problemet med FYROM : s namn , som , vilket ni säkerligen känner till , är föremål för en tvist med Grekland och för förhandlingar mellan de två länderna sedan mer än fyra år tillbaka , under FN : s generalsekreterares beskydd och inom ramen för säkerhetsrådets relevanta resolutioner , men även för ett kontraktsåtagande från parternas sida , på grundval av artikel 5 i det så kallade interimsavtalet från 1995 .
Jag anser det dock vara på sin plats att säga att den europeiska sidan , med anledning av de kommande förhandlingarna och slutandet av associeringsavtalet , för regeringen i Skopje bör betona nödvändigheten av att denna visar upp den lämpliga , konstruktiva politiska viljan och konstruktivt bidrar till att samtalen i New York slutförs på ett framgångsrikt sätt .
Jag vill hoppas att en sådan europeisk begäran , framförd parallellt med att man förklarar de svårigheter som ett eventuellt fortsatt dödläge kan leda till med avseende på slutförandet och tillämpningen av associeringsavtalet , kommer att ges erforderlig uppmärksamhet och utvärderas på lämpligt sätt av regeringen i Skopje , så att denna på motsvarande sätt svarar mot , å ena sidan , den tillmötesgående hållning som Grekland har uppvisat i frågan och , å andra sidan , mot den allmänt uttalade föresatsen och viljan hos alla Europeiska unionens medlemmar , inklusive Grekland , att underlätta och underbygga FYROM : s väg mot det enade Europa .
För , herr talman , jag tror inte att det faktum att det faktiskt existerar väl fungerande dagliga förbindelser , kontakter och kommunikation mellan FYROM och Grekland , såväl på det bilaterala som det multilaterala planet , främst tack vare de praktiska bestämmelserna i interimsavtalet , jag tror inte , skulle jag vilja säga , att det räcker för att de villkor och kriterier på god grannsämja som krävs för bland annat förhandlingar om och slutande av associeringsavtalet skall anses vara uppfyllda .
Tvärtom tror jag att ett sådant krav kan anses vara uppfyllt först efter att en de jure fullständig normalisering av förbindelserna mellan FYROM och alla dess grannländer har ägt rum .
Någonting sådant , i kombination med en nödvändig förbättring av vissa delar av landets inrikespolitiska situation , på området för minoriteter och de demokratiska institutionerna , kommer att komplettera den bild av politisk mognad som FYROM faktiskt uppvisar i övrigt och som har gjort att en förstärkning av förbindelserna med vår europeiska familj är välkommen .
Herr talman !
I den form som Swoboda har analyserat det , tas i dag med det avtal som vi diskuterar i dag - och som vi skall , hoppas jag , rösta igenom i morgon - det andra politiskt positiva steget , efter stabilitetspakten för regionen .
Det har även tagits ett litet steg , som hör samman med det partiella upphävandet nyligen av embargot mot Jugoslavien , vilket beslutades av våra 15 regeringar .
Mina damer och herrar , kolleger !
Regionen har befunnit sig i upplösning i ungefär tio år .
De tio åren , oavsett om man ser på dem som historisk eller som politisk tid , är en mycket lång tid .
Under dessa omständigheter är det alltså ett misslyckande i sak .
I den meningen är det avtal som vi skall rösta om i morgon och som faktiskt kommer att bidra till stabiliteten i regionen följaktligen ett steg i rätt riktning .
Före detta jugoslaviska republiken Makedonien ( FYROM ) är i själva verket en miniatyr av det tidigare Jugoslavien .
Oberoende av var den ena eller den andra minoriteten dominerar .
Ur den synvinkeln är det faktum att republiken fram till i dag har stått emot all påverkan från den omgivande miljön någonting mycket positivt , och inte under några omständigheter får någon av oss , någon stat , någon politik , någon åsikt - i ett försök att lösa andra problem - driva denna lilla demokrati till inre splittring , denna lilla demokrati som - vilket måste betonas - har institutioner som den kan utveckla ytterligare och därigenom bli en verklig demokrati .
I regionen har det till och från funnits flera typer av politiska modeller , och Europeiska unionen måste vara vaksam så att den inte - av ren tanklöshet - bidrar till att det byggs bananrepubliker på andra platser .
Vi måste veta att vi när vi söker allierade i denna region inte varje gång måste välja bland de som erbjuder sig .
Vi måste välja de som är moderata , som är vidsynta , som vill se fred och stabilitet i regionen .
Jag hoppas och önskar och är nu säker på att Europeiska unionen , med mognad och med de åtgärder som den har börjat vidta , sakta , sakta kommer att bygga upp den nödvändiga miljö som unionen själv behöver i hela regionen .
Vi får inte lura oss själva ; ett Europa med en region som är underutvecklad på grund av spänningar , på grund av olika missuppfattningar , på grund av motsättningar , på grund av konflikter mellan etniska grupper kommer under inga omständigheter att vara ett Europa som på sitt territorium har uppnått en nivå som kontinenten själv är nöjd med .
Hur som helst vill jag - nu i egenskap av grek - informera vissa kolleger som jag har lyssnat till om att många av talen rör sig i andra tider och på andra platser .
I dessa har man inte alls tagit hänsyn till de nya omständigheter som har formats i regionen , de nya positiva omständigheterna .
Vilket i väldigt många fall har skett efter initiativ av Grekland .
Och ni bör veta att det land som samarbetar mest av alla med den före detta jugoslaviska republiken Makedonien , det land i regionen som har de bästa förbindelserna med den före detta jugoslaviska republiken Makedonien är Grekland , och det har i mycket hög grad bidragit till stabiliteten i regionen .
Jag säger detta helt enkelt för att vi skall veta hur situationen ser ut i dag .
Herr talman !
Souladakis redogörelser tycks mig mycket förnuftigare än andra kollegers redogörelser från samma medlemsstat .
Låt mig säga i klartext att den som försöker göra överenskommelsen med Makedonien beroende av en lösning på namnfrågan i sin egen anda inte bara har Makedonien mot sig , utan även alla andra medlemsstater i Europeiska unionen .
Jag vill också vara tydlig och säga att han därmed skadar sitt eget lands intressen mycket svårt .
Det ligger i vårt intresse att det blir en stabil fredsordning på Balkan , och vi har chanserna , även om stabilitetspakten hotar att förvandlas till ett lik som aldrig har levat .
Jag hoppas att så inte blir fallet , men risken finns .
Just därför är det absolut nödvändigt att vi , EU , går bilateralt till väga med de enskilda staterna och att vi ger Makedonien ett tydligt europeiskt perspektiv .
Därför hälsar jag Swobodas utmärkta betänkande och i synnerhet punkt 12 i betänkandet som helt klart visar upp ett europeiskt , ett EU-perspektiv för Makedonien .
Jag anser att detta är viktigt , det måste ske , utan att för den skull hemfalla åt illusionism .
Vi vet att detta inte går från en dag till en annan , men att tydligt säga att Makedonien är ett otvetydigt europeiskt land och därmed har rätt att vara medlem i Europeiska unionen är en mycket viktig förtroendeskapande åtgärd .
Jag anser att vi har en enastående chans att stärka en demokrati som inte bara har fått till stånd en för detta område unik multietnisk regering , utan som även utvidgar det kommunala självstyret , reformerar rättsväsendet och näringslivet , och det under de svåraste villkor efter nationalism , kommunism och krig .
Jag hade äran att för några år sedan bjuda hit den nuvarande statschefen och den nuvarande ministerpresidenten som privatpersoner .
De hade då fortfarande stora problem med att bygga upp sina olika kontakter här .
Jag är mycket lycklig över att de har hållit vad de då lovade : att bygga upp en i grunden europeisk demokrati .
Vi måste tacka dem för att de i en mycket kritisk tid förra året som sagt spelade denna viktiga roll vid en strategiskt avgörande punkt vad gäller fred , stabilitet och demokrati .
Därför är vi inte bara de som ger , utan vi har också tagit , och vi är skyldiga makedonierna ett tack för att de då utförde ett avgörande europeiskt uppdrag .
Därför är det viktigt att avtalet förhandlas och ratificeras snabbt , att EU : s informationscentrum , den officiella delegationen , öppnas snabbt , att vår kommissionär enligt vad jag hör snart reser dit samt att vi öppnar upp ett entydigt europeiskt perspektiv åt detta land , liksom Swobodabetänkandet gör . .
( EN ) Det har varit en mycket intressant allmän debatt om Balkan som helhet .
Den blev inte sämre för det , men jag hoppas att ni förlåter mig för att jag i mycket hög grad koncentrerar mig på betänkandet , eftersom det finns några ytterst viktiga frågor som jag vill beröra .
Det gläder mig mycket att kunna framföra kommissionens synpunkter om betänkandet .
Det är ett mycket användbart betänkande .
Det är ett enastående bidrag från Swoboda och hans kolleger .
Vi är mycket tacksamma för hans engagemang i denna fråga , liksom för det engagemang som har visats av vissa av hans kolleger , av vilka några är här i kammaren i kväll - Pack , Lagendijk med flera .
Jag är mycket nöjd över att våra övergripande förbindelser med " FYROM " är så goda .
Jag hoppas att Dupuis - både han och hans tolk - förlåter mig för att jag använder termen i en anda av hjärtligt samförstånd .
Europeiska unionens förträffliga företrädare i landet har bidragit till detta .
Han har varit en pålitlig vän för parlamentet och till stor nytta för kommissionen .
Den nära förestående starten för förhandlingarna om ett stabiliserings- och associeringsavtal är det tydligaste exemplet på våra goda förbindelser .
Ett annat bra exempel är den före detta jugoslaviska republiken Makedoniens ( FYROM ) samarbete i återuppbyggnaden av Kosovo .
Jag är tacksam mot myndigheterna i Makedonien för deras hjälp under de senaste veckorna med att klara av de betydande svårigheterna med kraftförsörjningen i Kosovo .
I likhet med de ärade ledamöterna , inser jag den stabiliserande roll som detta land har spelat under tragedin på Balkan , särskilt när det gäller integreringen av den albanska minoriteten i landets politiska och sociala liv .
Jag träffade den nyvalda presidenten , Georgievski , för några veckor sedan , och jag blev - liksom andra har blivit - oerhört imponerad av hans engagemang för ett multietniskt och pluralistiskt samhälle .
Låt mig berätta var vi står i dag i dessa förhandlingar , som andra länder - vilket Lagendijk sade - i regionen följer med stort intresse .
Den 24 januari i år antog rådet sina förhandlingsdirektiv för ett stabiliserings- och associeringsavtal med före detta jugoslaviska republiken Makedonien .
Detta utgör det viktigaste steget framåt i den stabiliserings- och associeringsprocess för västra Balkan som kommissionen startade i maj 1999 .
Låt mig klargöra huvudpunkterna i dessa förslag till direktiv .
De omfattar inbegripandet i avtalet av åtgärder för att upprätta en politisk dialog med FYROM .
De omfattar bestämmelser för ökat regionalt samarbete , inklusive utsikten att upprätta frihandelsområden mellan länderna i regionen , fast jag måste göra det tydligt och klart att det inte är fråga om något försök att återskapa staten Jugoslavien .
De omfattar utsikten att upprätta ett frihandelsområde mellan Europeiska unionen och dem inom en tioårsperiod från det att avtalet träder i kraft .
De omfattar bestämmelser om rörlighet för arbetstagare , etableringsfrihet , tillhandahållande av tjänster , löpande betalningar och rörlighet för kapital .
De omfattar ett åtagande av FYROM att tillnärma landets lagstiftning till Europeiska gemenskapens lagstiftning , i synnerhet på vissa av den inre marknadens nyckelområden , och de omfattar bestämmelser om samarbete med FYROM på en stor mängd områden , inklusive rättsliga frågor och inrikesfrågor .
I kommissionen gör vi nu de nödvändiga förberedelserna , så att förhandlingarna kan påbörjas i mars .
Jag skall besöka FYROM den andra veckan i mars .
Jag hoppas kunna sätta processen i rörelse då , även om de formella förhandlingarna kommer att starta mycket kort därefter .
Under detta besök kommer jag också att uppgradera vår representation i FYROM , någonting som har rekommenderats av ärade ledamöter och andra .
Vårt riktdatum för att slutföra förhandlingarna är december i år , men detta kommer i mycket stor utsträckning att vara beroende av förhandlarnas goda vilja och beslutsamhet .
Avtalet skulle kunna träda i kraft om tre till fyra år räknat från i dag med hänsyn till den som krävs för ratificering i medlemsstaternas parlament .
Jag skulle helt kort vilja kommentera ett antal andra punkter i resolutionsförslaget .
Vi accepterar att avtalet i en viss utsträckning bör tjäna som ett exempel för andra , liknande avtal , även om vi självklart också måste ta hänsyn till det faktum att vi har att göra med olika länder , som vart och ett har sin egen identitet och sina egna angelägenheter .
Jag delar den allmänt spridda åsikten att vi bör behandla varje land efter deras meriter i stället för att binda upp alla till det långsammaste landets takt då det gäller utvecklingen av förbindelserna med unionen .
Det har aldrig varit avsikten .
Själva det faktum att förhandlingarna först startar med FYROM , före de andra länderna , är ett bevis på att vi kan göra - och att vi gör - åtskillnad .
Angående den bestämmelse om regionalt bistånd som hänvisas till i betänkandet , håller vi med om att vår tekniska och ekonomiska hjälp till en del bör gå till projekt med en gränsöverskridande eller regional dimension .
Vi håller med om att det bör finnas en utvecklingsklausul om utsikten till EU-medlemskap i stabiliserings- och associeringsavtalet .
Det skulle spegla Europeiska unionens syn på dess förbindelser med länderna på västra Balkan , såsom den formuleras i slutsatserna från Europeiska rådets möte i Köln .
Vi instämmer fullständigt i behovet av att decentralisera våra hjälpprogram i största möjliga utsträckning .
Vad beträffar uppgörelserna som omfattar Europeiska unionens hjälp till västra Balkan , tror jag att ledamöterna känner till att vi håller på att utarbeta en ny förordning , för att förenkla och strömlinjeforma programmens förvaltning och för att få in allting under en förordning .
Jag är medveten om att det finns en oro i FYROM och på annat håll över att Phare-programmet upphör i dessa länder och , framför allt , över att anknytningen till namnet Phare går förlorad .
Jag noterar med betydande oro vad ledamöterna säger i fråga om detta .
Jag skall se över frågan en gång till , fastän jag bör påpeka att det medför en risk för verklig förvirring att ha två Phare-program i gång samtidigt .
Jag vill emellertid betona att oavsett vad programmet kallas , är vårt åtagande att integrera FYROM och dess grannar i den europeiska familjen starkare än någonsin .
Rent allmänt är jag övertygad om att ledamöterna i denna kammare delar min belåtenhet över att Makedonien har nått detta stadium relativt snabbt .
Jag hoppas att de andra länderna i regionen kommer att fördubbla sina ansträngningar för att göra liknande framsteg .
Jag ser fram emot många liknande debatter om detta under de närmaste åren , vilka , hoppas jag , skall präglas av framgång för det som vi försöker göra på Balkan , som , i mina ögon , förblir det viktigaste avgörande provet på vad Europa kan åstadkomma på sin egen tröskel .
( Applåder ) Tack så mycket , kommissionär Patten .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Avtal om kommittéförfarandet Nästa punkt på föredragningslistan är betänkande ( A5-0021 / 2000 ) av Frassoni för utskottet för konstitutionella frågor om överenskommelsen mellan Europaparlamentet och kommissionen om de förfaranden som skall tillämpas för rådets beslut av den 28 juni 1999 - " kommittéförfarandet " ( 1999 / 468 / EG ) . .
( IT ) Herr talman !
I och med att vi godkänner detta avtal med kommissionen om hur rådets beslut om kommittéförfarandet skall tillämpas , avslutas ett ärende som under cirka två år har följt parlamentet och ett antal personer med ett passionerat intresse för denna fråga , personer som är utspridda inom unionens olika institutioner och som vissa inte skulle tveka att kalla masochister .
Ända sedan 1993 har sätten att utöva de olika behörigheter som delegeras av kommissionen , och framför allt den mystiska och kanske till och med suspekta verksamhet som kallas kommittéförfarandet , lett till konflikter och misstro mellan de olika institutionerna , något som riskerade att få allvarliga konsekvenser för lagstiftningsprocessen .
Det är av den anledningen som , i enlighet med förklaring nr 31 som bilagts Amsterdamfördraget , unionens institutioner har inlett ett komplicerat förhandlings- och samrådsarbete som utmynnat i rådets beslut att revidera det gamla systemet på ett ganska grundligt sätt , även om det för oss inte alls är helt tillfredsställande .
Framför allt omfattar beslutet ett förslag om att parlamentet skall ha vissa kontrollmöjligheter , dvs. man skall kunna slå larm om en åtgärd som genomförs till följd av en rättsakt som godkänts genom medbeslutande skulle kränka den beslutanderätt som delegerats till kommissionen .
Under den långvariga förhandlingen mellan institutionerna - där parlamentet har deltagit aktivt tack vare föredragandens , Adelaide Agliettas , arbete - var det underförstått att Europaparlamentet och kommissionen skulle sluta ett interinstitutionellt avtal om hur vissa aspekter av det nya beslutet skulle tillämpas .
Och detta skulle ske , å ena sidan , för att förtydliga vissa frågor som rådet inte hade för avsikt att åter ta upp i beslutet och , å den andra , för att på ett närmare sätt organisera informations- och kontrollsystemet när det gäller hur åtgärderna genomförs .
Under trepartssamtalen den 6 oktober 1999 i Strasbourg godkände Europaparlamentets talman och kommissionens ordförande idén att snabbt sluta ett sådant avtal .
Vi anser att vi har respekterat det åtagandet , som för övrigt har underlättats av det klimat av förtroende och ömsesidig respekt som kännetecknat samtliga förhandlingar med kommissionen .
De frågor som tas upp i avtalet är i huvudsak två : å ena sidan informationen till Europaparlamentet , ett conditio sine qua non för att parlamentet verkligen skall kunna utöva sin interventionsrätt i enlighet med artikel 8 i beslutet .
Den informationen har hittills getts i form av pappersdokument som skickats på ett osystematiskt vis , och många gånger på parlamentets eget ansvar , och informationen har varit oanvändbar för våra tjänstemän .
Från och med nu kommer informationen att lämnas via ett elektroniskt system som kallas Circa , som Europaparlamentet kommer att ha tillgång till och som kommer att innebära en verklig revolution , inte bara för oss , utan även - det är jag övertygad om - för kommissionen .
Å andra sidan preciserar artikel 8 i rådets beslut vare sig hur eller när Europaparlamentet skall slå larm , dvs. utöva sin begränsade kontrollmakt .
I artiklarna 6 och 7 i avtalet föreskrivs att Europaparlamentet i princip skall godkänna en resolution som motiverats i plenarsammanträde och att parlamentet har en månad på sig för att utnyttja sin rätt att ingripa innan kommissionens förslag till åtgärder godkänns .
Men det är inte alltid möjligt att vänta en månad innan en regel skall börja tillämpas , detta är vi alla medvetna om .
I avtalet ingår därför också en klausul om brådskande förfarande , som ger det ansvariga utskottet en möjlighet att ingripa .
Låt mig avslutningsvis understryka att för att bedöma om detta är ett bra avtal eller inte , så måste vi vänta och se hur det fungerar i verkligheten .
Europaparlamentet borde skaffa resurser , som man för närvarande inte förfogar över , för att garantera en effektiv uppföljning av verkställandet och en effektiv kontroll , och kommissionen borde acceptera att omorganisera vissa av sina rutiner för att garantera parlamentet en effektiv kontroll och en användbar information .
Slutligen kan det vara lämpligt att påminna om att under alla förhållanden så är för Europaparlamentets del den verkliga lösningen på problemen med kommittéförfarandet att ändra det förfarande för hur reglerna skall genomföras som anges i fördragen , samt en progressiv avveckling av kommittéerna , vilkas existens utgör en anomali som starkt begränsar kommissionens verkställande makt och som kan äventyra Europaparlamentets makt när det gäller lagstiftningsarbetet .
Herr talman , kära kolleger !
Kommittologi är ett begrepp som inte säger de flesta människor någonting , och endast fåtalet vet vad det innebär .
Det för tankarna till hemliga förbund och konspirationer , och så var det också förr .
Dock döljer sig bakom begreppet ingenting annat än fastställandet av villkoren för tillämpningen av de genomförandebefogenheter som anförtrotts kommissionen .
Villkoren för dessa genomförandebefogenheter består i ett begränsat antal kommittéförfaranden .
Fram till Amsterdamfördraget fanns det cirka 20 varianter av dessa kommittéförfaranden , vilket varken bidrog till klarhet i tillämpningen av lagstiftningen eller till genomsynlighet för medborgarna .
Tvärtom , under en lång tid blev inte ens självaste Europaparlamentet informerat .
Det första framsteget i kampen för mer öppenhet i denna kommittédjungel bestod för Europaparlamentets del i att man nu åtminstone informeras om allt det som Europeiska kommissionen har för avsikt att reglera inom ramen för dessa olika kommittéer .
Detta skedde genom brevväxlingen mellan Plumb och Delors 1988 .
Ett ytterligare steg i riktning mot öppenhet och delaktighet för Europaparlamentet blev sedan det så kallade modus vivendi av den 20 september 1994 , där parlamentet inte bara beviljades rätt till information , utan också en viss möjlighet att inlägga protester .
Därmed fick parlamentet även kontrollmöjligheter .
Med Amsterdamfördraget har situationen förbättrats avsevärt såtillvida att antalet kommittéförfaranden - liksom Europaparlamentet länge hade krävt - begränsades drastiskt till tre förfaranden , nämligen förvaltningsförfarandet , det föreskrivande förfarandet och det rådgivande förfarandet .
De informations- och kontrollrättigheter som har beviljats Europaparlamentet tidigare måste nu efter Amsterdamfördraget på nytt fastställs skriftligt i ett interinstitutionellt avtal .
Vår föredragande Frassoni har gjort ett mycket noggrant arbete och visat på vilka frågor om detta interinstitutionella avtal som måste redas ut och vilka förvaltningsförfaranden inom parlamentet som eventuellt måste ändras .
Ett nyckelproblem är tidsfaktorn .
När parlamentet informeras måste parlamentet , när man önskar ta ställning , i regel göra detta inom en mycket kort tidsfrist på fyra veckor .
I frågor som rör hälsa och säkerhet för människorna i Europeiska unionen måste Europeiska kommissionen som fördragens väktare och den enda institution som innehar initiativrätten vara i stånd att reagera med mycket kort varsel , i nödfall inom ett fåtal timmar eller dagar .
Trots det måste vi värna om Europaparlamentets rätt till information och eventuell reaktion .
Föredraganden visar på mycket användbara lösningar på dessa problem , vilka jag och min grupp stöder helt .
Jag har nu bara en bön till .
I den tyska texten under punkt 2 kan översättningen missförstås , och jag ber eftertryckligen om att detta rättas till , även i efterhand av de personer som ansvarar för tryckningen .
Enligt min mening bör det i stället för " weitergeführt werden müssen " ( måste föras vidare ) heta " erhalten bleiben müssen " ( måste upprätthållas , bevaras ) .
Detta är inte tydligt i den tyska texten .
Jag ber om att detta ses över igen .
I övrigt tackar jag vår föredragande hjärtligt .
Det är ett svårt ämne , och jag hoppas att vi har sett till så att vi nu kan sköta det bättre .
Herr talman !
Jag gratulerar föredraganden till hennes betänkande .
Jag måste tillägga att det är en välkommen förändring att se Frassoni vara i en så försonlig sinnesstämning och villig att kompromissa med de andra institutionerna .
När det gäller regeringskonferensen , är hon en av de personer som fransmännen kallar " les pures et dures " : inga kompromisser , inga uppgörelser med de andra institutionerna ; vi skulle hellre se hela saken blockeras än att kompromissa om våra ståndpunkter .
Men ändå är hon här villig att acceptera de steg framåt som har gjorts , vilka är långt från parlamentets ursprungliga ståndpunkter i frågan om kommittéförfaranden .
Låt oss komma ihåg vad som står på spel i denna fråga .
Parlamentet hade fyra huvudsakliga invändningar mot kommittéförfarandesystemet i den form det hade före det nya rådsbeslut som kompletteras av det interinstitutionella avtalet .
För det första är hela systemet dunkelt .
Det är inte öppenhet när hundratals kommittéer sammanträder med hemliga föredragningslistor och när ingen vet vilka personer som ingår i kommittéerna .
Här görs det ett verkligt steg framåt med det nya systemet som man har enats om .
Vi skall få veta vilka personer som ingår i de olika kommittéerna .
Vi skall få veta när de sammanträder .
Vi skall få ta del av föredragningslistorna .
Vi skall få ta del av de handlingar som sänds till dem .
Hela systemet kommer att bli mer öppet och genomblickbart - låt vara fortfarande ganska komplicerat .
Så det är åtminstone ett steg framåt .
Vår andra invändning är att systemet var mycket restriktivt med avseende på kommissionen .
Vi antar lagstiftning i Europeiska unionen .
Vi förväntar oss att kommissionen skall genomföra den .
Men sedan har vi ett system som är utformat så att det hindrar kommissionen och gör det svårare - särskilt det som kallades " contre-filet " systemet , enligt vilket rådet kunde blockera kommissionen med en enkel majoritet , även då rådet inte kunde finna alternativ till den aktuella genomförandeåtgärden .
Även här har det åtminstone gjorts vissa framsteg .
Rådet kommer inte längre att kunna blockera genomförandeåtgärder på obestämd tid efter tremånadersperioden , såvida det inte har en kvalificerad majoritet för att blockera dem , med andra ord , såvida det inte finns ett betydande motstånd bland medlemsstaterna som är företrädda i rådet .
Det är ett förnuftigare system .
Även detta är ett steg framåt .
Men i fråga om våra två andra invändningar är vi inte lika nöjda .
Den första invändningen gäller det system med vilket kommissionen övervakas , granskas , kontrolleras , om ni så vill , av en enda kommitté som utnämnts av medlemsstaterna eller rådet , inte av parlamentet .
Den lagstiftande myndighetens två delar , rådet och parlamentet , borde vara jämlika .
Vi tilldelar kommissionen genomförandebefogenheter , men sedan är det bara ett av rådet eller medlemsstaterna utnämnt organ som kan blåsa i visselpipan och säga nej till kommissionen och stoppa genomförandeåtgärden .
Parlamentet har ingen motsvarande maktbefogenhet .
Det är sant att vi nu ges ett första frö till en sådan befogenhet med det nya systemet .
Vi skall erhålla alla de förslag till genomförandeåtgärder som vidarebefordras till en kommitté samtidigt som de sänds till kommittén .
Vi kommer att ha möjlighet att granska , debattera och ifrågasätta .
Men vi kommer endast att ha rättighet att formellt bestrida kommissionen om vi anser att den har överskridit det bemyndigande som vi har gett kommissionen i lagstiftningen .
Med andra ord kan vi bestrida åtgärden för att det medför att befogenheterna , men vi kan inte bestrida innehållet i åtgärden .
Och i en demokrati borde parlamentet kunna bestrida innehållet .
Inte för att det är någonting som vi gör varje vecka .
Vi strävar inte efter att fördjupa oss själva i genomförandebeslut , men det är en demokratisk säkerhetsanordning att vi skall kunna göra det vid de få tillfällen som det verkligen skulle vara nödvändigt .
Detta saknas i det nya systemet , eller så är det bara där i embryoform .
Avslutningsvis , vår fjärde invändning är att om en genomförandeåtgärd blockeras genom kommittéförfarandesystemet , återförvisas det , men inte till den lagstiftande myndighetens två grenar , utan enbart till rådet , som har rättighet att vidta en eventuell alternativ åtgärd .
Detta är inte riktigt .
Båda grenarna - rådet och parlamentet - antar den lagstiftning med vilken kommissionen tilldelas genomförandebefogenheter .
Om sådana genomförandeåtgärder återförvisas , bör det vara till båda grenarna , inte bara till den ena .
På det hela taget har vi ett system som har gått framåt .
De kompletterande aspekterna som härrör från den interinstitutionella avtalet med kommissionen är välkomna , men det kan inte ändra rådets grundläggande beslut .
Även här har vi frivilligt - eftersom det inte var någonting som skedde automatiskt - gett upp Plumb-Delors-avtalet som en del av den övergripande kompromissen .
Vi har gått med på att avstå från bestämmelserna i det .
Vi måste vara väldigt vaksamma på det som tidigare omfattades av det avtalet och som nu inte helt omfattas av det nya beslutet .
Vi måste vara mycket vaksamma .
Så det är ett steg framåt .
Min grupp accepterar det motvilligt som ett steg framåt .
Vi känner inte alls samma entusiasm för att kompromissa som Frassoni .
Vi inser att det finns begränsningar och att frågan utan tvekan kommer att komma tillbaka inom några få år .
Om vi vill ha en union som verkligen är demokratisk och öppen , måste vi ta upp detta ämne igen . . - ( ES ) Herr talman !
Jag vill börja med att tacka föredragande Frassoni för hennes insats .
Att arbeta med kommittéförfaranden är aldrig lätt .
Schleicher har hänvisat till den typ av magi som vi alltid har talat om , om kommittéerna .
Det stämmer att det alltid har varit en mycket invecklad process till följd av tidigare historiska beslut som man till slut måste rationalisera någon gång .
Enligt min uppfattning innebär den överenskommelse som kommissionen och parlamentet har kommit fram till en tydlig rationalisering av processen .
Vi anser att den tillgodoser parlamentets grundläggande intressen .
Corbett har tagit upp några orosmoment .
Han säger att vissa av dem har fått en lösning och andra inte .
Jag skulle nog vilja påstå att de kommissionen har kunnat lösa har fått en lösning .
Det som tas upp av Corbett är andra premisser som inte omfattas av rådets beslut , och där vi tyvärr inte kan gå längre .
I vilka avseenden har vi gjort framsteg ?
Utan tvekan i en grundläggande fråga som Frassoni har lyft fram , nämligen att vi har ett automatiskt informationssystem .
Detta automatiska informationssystem kommer att möjliggöra två aspekter som är av särskilt intresse för parlamentet .
Å ena sidan för att få information om hur kommittéerna har fungerat , deras sammansättning , dagordning , framställningar , osv . , och å andra sidan insyn angående konkreta beslut .
Jag anser att det är en bra överenskommelse .
En bra överenskommelse som utan tvivel ökar insynen i processen .
Från och med nu kommer saker och ting att gå lättare .
Den överenskommelse vi uppnår i dag bör emellertid inte betraktas som en steg bakåt vad beträffar avtalet om Delorsplanen .
Corbett tog upp frågan , men den nya modellen är mycket mer omfattande , annorlunda till följd av den nya situationen och i vårt tycke betydligt mer enhetlig .
Vi har redan påbörjat arbetet .
Låt oss hoppas att det leder till goda resultat .
Å andra sidan betraktar vi även andra framsteg som positiva .
Vi överträffar i vissa avseenden avtal som redan är föråldrade och vi försöker genom att återanpassa gamla förfaranden till den nya situationen att rensa bort sådant som finns kvar från förr .
Kommissionens slutsats är att det är en bra överenskommelse , som vi vill tacka de parlamentariker för - och då i synnerhet Frassoni - som har arbetat med denna .
Vi hoppas att man i det nya klimatet har lyckats uppnå det resultat man eftersträvade , nämligen en ökad öppenhet och större kännedom om de beslut kommissionen fattar i kraft av sina verkställande befogenheter .
Tack så mycket , kommissionär Solbes Mira .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Protokoll om förfarandet vid alltför stora underskott Nästa punkt på föredragningslistan är betänkande ( A5-0013 / 2000 ) av Knörr Borràs för utskottet för ekonomi och valutafrågor om förslaget till rådets om en ändring av förordning ( EG ) nr 3605 / 93 om tillämpningen av protokollet om förfarandet vid alltför stora underskott som är fogat till Fördraget om upprättandet av Europeiska gemenskapen ( KOM ( 1999 ) 444 - C5-0174 / 1999 - 1999 / 0196 ( CNS ) ) .
( ES ) Herr talman !
Jag har nöjet att även få hälsa på den spanske kommissionären Solbes som jag vid mer än ett tillfälle har gratulerat , både inom och utanför parlamentet , till hans utmärkta insats i konungariket Spanien vad gäller den europeiska konvergensen .
I förslaget till förordning om ändring av förordning ( EG ) nr 3605 / 93 om tillämpningen av protokollet om förfarandet vid alltför stora underskott som är fogat till Fördraget om upprättandet av Europeiska gemenskapen tas frågan upp om en anpassning till räkenskapssystemet ENS 95 vilket , som ni vet , kom att ersätta det tidigare Europeiska nationalräkenskapssystemet från 79 .
Förslaget inbegriper i synnerhet nya finansiella utgiftsområden , enhetlighet i beräkningen av kvoten mellan underskott i den offentliga sektorns finanser och BNI mot bakgrund av ENS 95 samt vikten av att ränteutgifter beaktas och av att dessa utgifter sinsemellan är jämförbara i enlighet med metodiken i ENS 95 .
Förslaget till förordning är , enligt min uppfattning , en aktualisering av definitionerna och en bedömning av somliga av de ekonomiska åtgärder som påverkar beräkningen av underskottet så som framgår av Maastrichtfördraget , där maximala procentsatser till marknadspriser för de offentliga förvaltningarnas underskott ställs i förhållande till bruttonationalinkomsten i unionens olika medlemsstater .
Hittills har staterna räknat ut BNI enligt metodiken i ENS 79 .
Den sista beräkning vi har tillgång till skedde i september 1999 och avsåg budgetåret 1998 .
Om föreliggande förordning antas kommer beräkningen i mars månad 2000 , den första beräkningen av underskottet för budgetåret 1999 , att ske med det nya systemet .
Man vet att medlemsstaterna- om man får uttrycka sig så - har skött sin uppgift , de har gjort en uppställning av sina nationella räkenskaper i enlighet med ENS 95 , och deras beräkningar har redan offentliggjorts .
Detta förfarande har inneburit att medlemsstaterna förutom att inbegripa en ny metodik även har genomfört en nominell revision av största delen av aggregaten och redovisningskalkylerna .
Denna revision är både ett resultat av att nämnda metodikändringar genomförts och att ett bättre statistiskt underlag tagits med i beräkningarna .
Dessa ändringar kan givetvis påverka medlemsstaternas statsfinanser vad beträffar den offentliga sektorns underskott .
Nu vill jag i all korthet tala om vilka de fem områden kan vara där de viktigaste ändringarna sker .
För det första , en anpassning av den definition av offentlig sektor som ingår i ENS 95 .
Detta är viktigt eftersom underskottet i den offentliga sektorns finanser beräknas på grundval av hela den offentliga sektorn .
Om man inte förfogar över de kriterier som är nödvändiga för definitionen av denna , kommer det att leda till avvikelser vid beräkningen av underskottet inom den offentliga sektorn i medlemsstaterna .
För det andra , underskottet - eller i förekommande fall överskottet - inom den offentliga sektorns finanser motsvarar den offentliga sektorns nettoupplåning eller finansiella sparande enligt definitionen i ENS 95 .
För det tredje , offentliga investeringar motsvarar den offentliga sektorns fasta bruttoinvesteringar enligt definitionen i ENS 95 .
För det fjärde , den offentliga sektorns skuldsättning och de flöden ( räntor ) som härrör från dessa skulder / tillgångar definieras i enlighet med ENS 95 .
Och slutligen för det femte , den aggregat som ligger till grund för beräkningen av underskottet skall vara bruttonationalinkomsten till löpande marknadspriser , uppskattad i enlighet med definitionerna i Europeiska nationalräkenskapssystemet 95 .
Kort sagt , kommissionens förslag visar enligt min uppfattning på en korrekt och konkret överensstämmelse mellan de kriterier som fastställs i Europeiska nationalräkenskapssystemet 95 som jag därför godkänner i sin helhet , precis så som det framlagts av kommissionen .
Herr talman , herr kommissionär , mina damer och herrar !
Låt mig säga direkt att min grupp välkomnar detta förslag eftersom den statistiska grunden för en ekonomisk och monetär union som koncentrera till stabilitet och reell tillväxt härigenom utformas mer harmoniserat , direkt jämförligt och mer exakt .
Vi har redan hört de olika områdena .
För mig är det avgörande att de statistiska uppgifterna från och med nu blir mer tillförlitliga och mer jämförliga .
Detta är nödvändigt därför att vi måste kunna lita på varandra : de olika organen inom Europeiska unionen och alla medlemsstater inom valutaunionen .
En anpassning av förfarandet är viktig av två anledningar .
För det första för den inre marknadens skull .
Tillförlitliga och direkt jämförbara data och statistik är rent allmänt av stor betydelse för en exakt skildring av situationen och utvecklingen på en inre marknad .
För det andra för den ekonomiska och monetära unionens skull .
Förordningen från 1993 som gäller tillämpningen av protokollet måste fås att harmoniera på nationell och regional nivå med metodiken för Europeiska nationalräkenskapssystemet .
Detta är oumbärligt för ett korrekt och tillförlitligt fastställande av underskotten .
Anpassningen kommer att göra det möjligt att åstadkomma en precis bedömning av underskotten och skuldnivån i medlemsstaterna .
Denna tekniska anpassning kommer att få mycket konkreta konsekvenser för staternas faktiska ställning eftersom siffrorna ändras automatiskt i förhållande till de offentliga underskotten .
Jag välkomnar även det faktum att deklarationen av underskotten för budgetåret 1999 som skall offentliggöras i mars 2000 redan utarbetas efter det nya Europeiska nationalräkenskapssystemet , vilket innebär att analysen baserar sig på ur ekonomisk synvinkel relevant , konsoliderat statistiskt material .
Men låt mig använda debatten även till att helt kort vädja till alla regeringar och politiska partier att göra allt för att förfarandet vid alltför stora underskott aldrig skall behöva tillämpas .
Det är bra att förfarandet finns .
Förfarandet är nödvändigt eftersom det skänker nödvändigt tyngd och trovärdighet åt våra villkor .
Medborgarna frågar : Vad händer om villkoren inte uppfylls ?
Med förfarandet och andra åtgärder kan vi bevisa att vi menar allvar med villkoren och med oss själva .
En andra väsentlig punkt gäller att vi måste satsa allt på att förhindra inte bara de alltför stora underskotten , utan offentliga underskott måste sänkas mer än så .
Jag vet vad jag talar om , och låt mig avslutningsvis säga varför jag är så glad över att vi för denna debatt !
I mitt eget land för vi för tillfället diskussioner om huruvida de upplysningar som förre finansministern har lämnat om underskottet motsvarar den faktiska verkligheten .
I mitt eget land , i Österrike , krävdes det 1995 ett nyval för att Maastrichtkriterierna skulle uppfyllas och den politiska partnern förmås att tänka om .
Jag måste också säga att år 2000 , då det ju talas så mycket om oss , misslyckades - jag säger tyvärr - koalitionsförhandlingarna med SPÖ ( Österrikiska socialdemokratiska partiet ) eftersom det besparings- och konsolideringsprogram som förhandlats fram bragdes på fall av det socialistiska partiet .
Inte minst var man tvungen att bilda den nya regeringen i Österrike därför att ÖVP ( Österrikiska folkpartiet ) vill fortsätta att garantera stabilitetskursen , därför att ÖVP vill fortsätta se till att Maastrichtkriterierna uppfylls liksom att de offentliga underskotten minskas , vilket vi här har kommit överens om .
Herr talman !
Det är bra om statistiska uppgifter inte bara är pålitliga , utan också är jämförbara .
Det är av stor betydelse , framför allt för det europeiska enandet och fullbordandet av den inre marknaden .
Därför är detta betänkande också ett politiskt laddat betänkande som vi vill framföra våra hjärtliga gratulationer till föredraganden för .
Det ger också anledning till ett par politiska kommentarer .
Stabilitetspakten är ett faktum i Europa .
Alla länder som deltar i euron har via denna stabilitetspakt förpliktigat sig att på medellång sikt sträva efter en budget som är i balans eller som uppvisar ett litet överskott .
Det skall naturligtvis inte innebära att det skulle kunna bli något mer eller något mindre om konjunkturen är något ogynnsam , men på lång och medellång sikt måste det handla om balans eller ett överskott .
Ju starkare de deltagande ländernas ställning blir , desto starkare kommer euron att bli .
Härigenom kommer treprocentsnormen sällan att överskridas , inte heller under konjunkturmässigt ogynnsamma omständigheter ; det är i alla fall så som resonemanget lyder .
Vi har alltid ansett att dessa kriterier måste vara strikt uppfyllda .
Det är av stor betydelse för att kunna göra EMU till en framgång även i framtiden .
Sträng efterlevnad av stabilitetspakten kan på så sätt bidra till att det uppstår en stablitetskultur i alla EMU-medlemsstater .
Vissa medlemsstater har vidtagit engångsåtgärder för att kunna uppfylla kriterierna .
Vi anser att medlemsstaternas budgetpolitik måste hållas under sträng tillsyn , så att åtgärderna hela tiden överensstämmer med andan i de ställda kriterierna .
Någon avmattning får inte tillåtas .
Vidare anser vi att ett minskat skattetryck och en minskning av statsskulden måste tillhöra prioriteringarna .
För det är ju så att vi fortfarande inte har upphört att övervältra bördorna på kommande generationer . .
( ES ) Herr talman !
Först av allt ett tack till föredraganden för hans fantastiska arbete .
Detta ämnesområde innehåller många facktermer och jag anser att Knörr har behandlat frågan med stor precision och ett stort yrkeskunnande .
Jag vågar inte försöka sammanfatta innehållet i vårt förslag bättre än han har gjort ; jag skulle endast vilja göra ett litet tillägg genom att säga att det förutom anpassningen till ENS 95 finns två mindre tekniska ändringar som Knörr känner väl till och som avser räntorna och skuldutvecklingen i utländsk valuta .
Det säger jag bara som en kommentar för att processen skall ses i sin helhet .
För det andra vill jag tacka Knörr för hans snabba insats .
Han har gjort ett mycket bra arbete på kort tid .
Det här är en viktig fråga , med tanke på de kommentarer som vi har fått .
Vårt syfte med den här bestämmelsen är inte att de statistiska uppgifterna skall bli trovärdiga och jämförbara - det är de redan - utan att de skall bli ännu mer trovärdiga och jämförbara .
Det är uppenbart att vi , tack vare att parlamentet har fattat beslut så snabbt , kommer att kunna beräkna siffrorna redan för mars månad med hjälp av de nya kriterierna .
Jag tror att slutresultatet kommer att bli bättre framöver .
Sifferuppgifterna kommer att vara mer tillförlitliga och jämförbara och jag tror att den oro som vissa av er har uttalat beträffande uppfyllandet av stabilitetspakten lättare kommer att kunna bedömas .
Denna förordning tjänar enbart som ett instrument .
Med hjälp av den kommer vi inte till kärnan av det problem precis som vissa av er har påpekat .
Däremot kan vi säga att vi har fått fram vilken problemets kärna är .
Stabilitetspakten existerar , låt oss nu fortsätta framåt genom att se till att de olika medlemsstaterna uppfyller den , även i en situation som den nuvarande , då resultaten är klart positiva i alla de medlemsstater där vi har undersökt situationen vad gäller stabiliteten i den offentliga sektorns underskott .
Däremot får vi inte sänka beredskapen .
Vi måste envist följa denna färdriktning som vi betraktar som grundläggande .
Än en gång , därför vill jag - och härmed avslutar jag mitt anförande - tacka för er hjälp så att vi kan mäta stabiliteten med en större fackmässig garanti och bättre möjligheter till jämförbarhet .
Tack så mycket , kommissionär Solbes Mira .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Euro : förstärkning av det straffrättsliga skyddet mot förfalskning Nästa punkt på föredragningslistan är betänkande ( A5-0020 / 2000 ) av Cederschiöld för utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor om förslaget till rådets rambeslut om förstärkning av det straffrättsliga skyddet mot förfalskning i samband med införandet av euron ( 5116 / 1999 - C5-0332 / 1999 - 1999 / 0821 ( CNS ) ) . .
Herr talman , kära fåtaliga , men desto mer välkomna kolleger !
Man kunde tro att det vid denna timma skulle vara ett oviktigt ärende som skall behandlas , men så är icke fallet .
Det är en handfast och konkret fråga .
Det handlar om vår gemensamma valuta .
Hur många här vet att den valutan förfalskas , och att vi har helt oacceptabla förhållanden ?
Vi kan inte tillåta att vår gemensamma valuta förlorar kraft genom att den förfalskas .
Därför har ECB , Ekofin , Europol , OLAF och kommissionären med ansvar för rättsliga frågor insett att det snabbt måste vidtas gemensamma motåtgärder för att fylla de luckor som lagstiftningen uppvisar .
Det är lätt att glömma att de gamla valutorna kan växlas in tjugo år efter det att den nya valutan har introducerats .
Därför är det viktigt att inkludera även dessa valutor i den straffrättsliga delen av detta åtgärdsprogram .
Det har parlamentet velat lägga till .
Rådet borde ha givit parlamentet den stipulerade tremånadersfristen även för det sista dokumentet som man tog fram i detta ärende , men vi är alla medvetna om hur brådskande det är att få dessa åtgärder i hamn .
Eftersom frågan skall beslutas om i mars i rådet , finns det anledning för parlamentet att nu ta ställning till förslaget , så att medlemsländerna hinner väga in även parlamentets ståndpunkter i det beslut som måste fattas i mars .
Om något land skulle börja krångla , drar det landet på sig ett ansvar för valutan som borde göra det landet ansvarigt , både moraliskt och ekonomiskt , om det skulle bidra till en försening .
Ett sådant agerande skulle medföra mycket badwill .
Den 1 januari 2002 är euron i omlopp .
Hela unionen måste ha samma skydd , ett skydd som förbjuder förfalskningar , inte endast av valutor i omlopp utan också av valutor som kommer att komma i omlopp .
Det är viktigt att i tid ha ett straffrättsligt skydd i alla länder som ser någorlunda likadant ut .
Kommissionen har föreslagit informationsåtgärder , förebyggande åtgärder , utbyte av erfarenheter och straffrättsliga åtgärder , som faktiskt innebär en viss nödvändig tillnärmning , nämligen att det lägsta acceptabla maxstraffet för valutaförfalskningar blir åtta år .
Även handel med falska valutor och innehav av förfalskningsutrustning kommer att kriminaliseras .
Vi får helt enkelt en miniminivå för det högsta straffet .
Eurons valörer är väl kända .
Modern datautrustning kan åstadkomma en hel del skada om vi inte skyddar oss .
Parlamentet har tillfört ett antal ändringsförslag till detta liggande förslag , bl.a. när det gäller domsrätt , som innebär att man endast får åtalas och dömas i ett land för samma brott .
Åtgärder mot företag som är inblandade i förfalskningar finns också med , vilket vi tillskyndar .
De nya kandidatländerna uppmanas också att anpassa sig till dessa regler .
Det har tagit två år för rådet och kommissionen att få fram detta förslag .
Det är absolut nödvändigt att beslutet nu tas i mars .
Att försena eller kanske till och med riskera skador på euron vore oförsvarligt .
Det vore också ett svek mot medborgarna som skall hantera de nya , obekanta sedlarna .
Särskilt tror man att falskmyntarna vänder sig mot länder som står utanför euron , där medvetenheten om den nya valutan är svagare .
Skyddsåtgärderna omfattar även dessa länder , och synpunkterna från dessa länder har fått väga tungt .
Därför kan man beteckna detta förslag som solidariskt och ömsesidigt i sitt ansvarstagande för olika intressen , vilket förpliktigar .
Rådet måste nu i mars möta upp och fatta detta beslut .
Tack kollegor för att ni lyssnade .
Tack även till dem som har bidragit till en snabb hantering i frågan ; jag tänker särskilt på PSE-gruppen .
Herr talman , ärade kollegor !
Jag vill börja med att tacka föredragande Charlotte Cederschiöld för ett bra betänkande , en utmärkt utgångspunkt för en förstärkning av det straffrättsliga skyddet mot valutaförfalskning inför eurons införande .
Euron sätts i omlopp den 1 januari 2002 och blir en av de viktigare valutorna i världens valutareserv .
På grund av dess betydelse på det internationella planet kommer euron att vara särskilt utsatt för förfalskning och plagiat .
Med det här förslaget till beslut kommer ett minimum av regler att fastställas genom att man försöker harmonisera straffrätten på området och förenkla och effektivisera tillämpningen för varje medlemsland .
Man räknar fortfarande med att skyddet för euron skall vara klart innan den sätts i omlopp , vilket för många länder kommer att täcka en lucka i lagen .
Jag vill uttryckligen stödja föredraganden i det hon säger om nödvändigheten av att utsträcka skyddet till att gälla även de nationella valutor som man kan fortsätta att växla in efter att de dragits tillbaka .
Varje stat måste därmed se till att effektiva straffpåföljder införs , påföljder som skall vara lämpliga och avskräckande för de brott som förutses i förslaget till rambeslut .
Beträffande förslaget om en maximigräns på åtta år för frihetsberövande straff , utgör detta enligt min mening inga som helst problem för mitt land som , trots att man i sin brottsbalk håller på att sänka det maximala straffet till fem års fängelse för valutaförfalskning , visade sig vara beredd att ta itu med respektive ändringsförslag .
Å andra sidan vill jag uppmana de få medlemsländer som fortfarande har vissa reservationer att lösa detta , så att vi snarast kan fatta ett beslut , precis som föredraganden vädjade om och av samma skäl .
Herr talman , med detta förslag till rambeslut har vi för första gången lagt fram ett gemensamt straffrättsligt förslag med lagar som skall tillämpas av de femton medlemsländerna samtidigt .
Därmed tar vi ett steg mot vårt mål att utveckla och konkretisera Europeiska unionen när det gäller området frihet , säkerhet och rättvisa , vilket också beaktades i Tammerfors .
Herr talman , ärade kolleger !
Jag behöver inte upprepa vad föredraganden har sagt , inte heller vad Coelho redan har redogjort för .
Allt är nämligen rätt och riktigt .
Euron kan lätt förfalskas .
Vi befinner oss i en riskabel övergångsfas där det straffrättsligt uppträder ett - jag antar i penningväsendets historia - väl unikt fenomen , nämligen att en valuta som ännu inte är tillgänglig , som ännu inte är i omlopp utan endast existerar som giromedel ändå redan kan förfalskas , men att valutaförfalskningen i nuläget ännu inte kan bestraffas på grund av just det faktum att valutan ännu inte är i omlopp .
Ett rätt komplicerat problem .
Det vill säga , man kan , om vi inte agerar snabbt - det har Cederschiöld rätt i - redan nu tillverka ett par falska euro och eventuellt slippa att ställas till svars för att dessa sätts i omlopp .
För en och annan , det tillåter jag mig att säga i förbigående , lär detta kunna vara en attraktiv chans .
Vad gör nu Europeiska unionen för att förhindra detta ?
En rad korrekta åtgärder , vilka Cederschiöld har beskrivit , men parlamentet behöver inte säga så mycket om innehållet i de rambeslut som Cederschiöld har beskrivit , inte så mycket om det betänkande hon har författat som om de förfaranden som tillämpas .
Europaparlamentet har av rådet , den absolut mest odemokratiska institutionen i Europa , rådfrågats på ett sätt som är ett hån mot begreppet demokrati .
Vi har fått en text översänd för samråd som rådet självt har knåpat på under en mycket lång tid , för övrigt endast till viss del med framgång - jag skall strax återkomma till detta .
Nu skall Europaparlamentet på tre månader ta ställning till detta komplexa , svåra , delvis motsägelsefulla dokument från rådet .
Det är endast tack vare kollegan Cederschiölds enorma insats liksom att Europaparlamentet avstår från att utnyttja sin demokratiska rätt att få tillräcklig tid på sig samt tillgång till alla texter på alla språk för att genomföra ett samrådsförfarande som vi nu kan få ett ställningstagande inom de tidsramar som rådet önskar och därmed komma fram till det beslut som skall fattas i mars .
I en så viktig fråga som valutaförfalskning , eller skyddet mot valutaförfalskning , och den straffrättsliga standardisering som det kräver , kan man egentligen inte arbeta i ett så svinaktigt tempo som rådet kräver att vi skall göra .
Därför vill jag nu på min grupps vägnar säga rent ut : Vi har diskuterat länge med kollegan Cederschiöld huruvida det kan vara vettigt att arbeta så här .
Vi har kommit fram till att så inte är fallet , men med tanke på hur viktigt ämnet är har vi ändå enats om att acceptera förfarandet .
Det råder ingen tvekan om att föreliggande rambeslut är ett steg framåt .
Det är bara det att den rättssäkerhet , som det egentligen var rådet som önskade - det har Cederschiöld redan utvecklat - inte kommer att uppnås helt i alla fall , för när det gäller den eftersträvade miniminivån , det lägsta godtagbara maximistraffet , och framför allt tillämpningen av en identisk straffrättslig norm i alla medlemsstater - även i de länder där euron ännu inte har införts men där den teoretiskt sett skulle kunna förfalskas - har bristerna inte avhjälpts .
Bland annat har de inte avhjälpts därför att rådet som vanligt inte kan handla mot sin egen natur utan även vid detta rambeslut föredrar att framhärda på regeringssamarbetsnivå när det gäller just det rättsliga samarbetet .
Därför är detta rambeslut - det skall jag gärna citera - också bara en komplettering till ett internationellt avtal som har 71 urvattnade år på nacken , nämligen avtalet av den 20 april 1929 om bekämpning av falskmynteri och därtill hörande protokoll .
Det här betyder att vad vi nu utarbetar som juridiskt underlag för att skydda euron inte görs där detta egentligen borde göras , nämligen på gemenskapslagstiftningens område , utan det görs som en komplettering till internationella överenskommelser som är 71 år gamla .
Huruvida detta kan vara Europeiska unionens framtid , framtiden för det rättsliga samarbetet i Europeiska unionen , det överlåter jag åt närvarande församling att avgöra .
Jag tackar för den uppmärksamhet jag har fått för vårt gemensamma nattliga program .
Herr talman !
Eurons införande skulle mycket väl ha kunnat vara en välsignad period för falskmyntare .
Medborgarna kommer i ett slag att förlora alla sina penningreferenser och riskerar därmed att lätt acceptera falska euro , då de ännu inte har lärt känna de nya så väl .
Det är således naturligt att rådet oroar sig över detta och söker föreskriva påföljder , i synnerhet straffrättsliga , för den här typen av brott , vilka skall kunna tillämpas i hela Europa .
För det ändamålet hade det utan tvekan kunnat nöja sig med en enkel resolution , där man rekommenderar medlemsländerna att anta nationella lagar med den innebörden .
Det är vad jag personligen hade trott var att föredra .
Men rådet - utan tvivel för att det saknar förtroende för vissa medlemmars nit - föredrog i stället att etablera ett mer tvingande rättsligt instrument på EU-nivå , dvs. ett rambeslut .
Och det är där svårigheterna börjar , eftersom straffrätten lyder under den nationella suveräniteten och eftersom Maastrichtfördraget inte föreskriver något specifikt för euron i det här sammanhanget , för att man inte ville skrämma väljarna genom att lasta båten för tungt .
Det utkast till rambeslut som presenteras för oss i dag försöker således dölja denna lucka genom att hänvisa till artiklarna 31 e och 34.2 b i fördraget .
Men dessa hänvisningar förefaller otillräckliga .
Artikel 31 föreskriver endast gemensamma minimiregler för straffrättsliga brott i ett begränsat antal uppräknade fall : organiserad brottslighet , terrorism och narkotikasmuggling .
Falskmyntning ingår inte .
Artikel 34 , ett resultat av Amsterdamfördraget , definierar endast den nya formen för rambeslut , men den tillämpas självklart bara på de befogenheter som unionen redan har .
Vi kommer därmed tillbaka till det tidigare nämnda problemet .
Med andra ord har rådet inte lyckats ge denna text en trovärdig rättslig grund .
Det är på något sätt ett försenat straff för den brist på ärlighet som rådet uppvisade då det presenterade Maastrichtfördraget för väljarna .
Jag skulle också vilja framhålla en mer allmän tanke .
För en tid sedan fick vi nästan under alla sammanträdesperioder behandla ett eller flera betänkanden om principfrågor kring euron .
Men sedan ett år tillbaka : inga alls .
Endast några mindre tekniska betänkanden , såsom det om förfalskningar .
Kommissionens meddelande om strategiska målsättningar för 2000-2005 , vilket vi debatterade i veckan , innehöll absolut ingenting om detta stora ämne , bortsett från en erinran , med en rad , om att mynten och sedlarna i euro kommer att sättas i omlopp den 1 januari 2002 .
Det är verkligen mycket tunt .
Ändå finns det många grundläggande problem som inte är lösta .
Vi kan till exempel nämna det oroväckande ointresset från allmänhetens sida ; att de penningpolitiska målen har reducerats till att endast omfatta inflationsbekämpning ; att man märkligt nog har upprättat en monetär federalism utan vare sig en finansiell eller skattemässig federalism ; de aktuella kandidatländernas status visavi euroområdet då de kommer att ha blivit medlemmar ; de internationella marknadernas villrådighet inför en valuta utan ett homogent befolkningsunderlag , osv .
Behöver man också erinra om att de investerare som har sålt dollar för att köpa euro har förlorat 20 procent sedan den 1 januari 1999 , 40 procent om de köpte obligationer och till och med 55 procent om de sålde yen för att köpa euro .
För dessa stackars investerare , herr talman , är även riktiga euro falska pengar .
Det är gigantiska problem , men här tycks de vara tabubelagda .
Jag vill gärna ta upp tråden från föregående talare .
Det finns några principfrågor som tränger sig på , därför att utgångspunkten är ju att den straffrättsliga regleringen är en nationell angelägenhet .
Straffrätten tillhör det enskilda samhällets kulturella tradition , och det är mycket svårt att komma fram till gemensamma definitioner av vad som avses med dessa juridiska grundbegrepp .
Jag uppskattar Cederschiölds arbete och jag utgår från hennes efterlysning - i samband med toppmötet i Tammerfors - av gemensamma definitioner och bestämmelser för vad som är straffbart , och vilka gemensamma sanktioner som kan komma ifråga .
Hon vill gärna utarbeta dessa sanktioner gemensamt för att komma fram till ett samstämmigt system för överträdelser som är särskilt relevanta för EU .
Men problemet är att det inte finns stöd för det - och detta har goda skäl , eftersom den straffrättsliga regleringen tillhör den nationella behörigheten .
I detta sammanhang vill jag ställa följande frågor till kommissionens och rådets företrädare : Är den rättsliga grund som åberopas tillräcklig ?
Enligt min uppfattning strider den helt klart mot och går långt utöver artikel 34.2 b , där rättsstödet fastställs för s.k. rambeslut , som är bindande för medlemsstaterna vad gäller de åsyftade målen , men där det överlåts till de nationella myndigheterna att bestämma form och medel för genomförandet .
Det som är karakteristiskt för det föreliggande förslaget till rambeslut är ju att man i detalj fastställer medlemsstaternas förpliktelser - det finns inte någon valfrihet när det gäller medlen och genomförandet .
Och enligt min uppfattning går detta utöver ramarna för stödet .
Jag vill gärna ha ett svar från kommissionen och rådet , därför att jag anser det vara uppenbart att det inte finns stöd i artikel 31 .
Herr talman , fru kommissionär !
Jag vill inleda med att hjärtligt gratulera och tacka föredraganden och även peka på att hon i sitt betänkande ju inte bara välkomnar förslaget till rambeslut , utan att hon också har föreslagit vissa ändringar som skall komplettera och förbättra texten , vissa ändringar som även har tagits upp av de olika talarna men som vi inte kan genomföra alla nu .
Hur som helst handlar det om att fortsätta historieskrivningen om eurons framgångar , och vi måste göra allt för att denna framgångsrika historia inte skadas eller ifrågasätts på grund av för svaga motåtgärder mot förfalskning - några första ansatser känner vi redan till .
Vi har alla pekat på att omställningsfasen också innebär osäkerhet och risker .
Därför måste också den planerade informationskampanjen som vi måste ägna oss mycket intensivt åt naturligtvis komma att spela en viktig roll vid sidan av arbetet mot förfalskningar , mot en vederbörlig tillämpning av bestämmelserna .
Men det gäller också frågor om samarbetet .
Vi behöver definiera den exakta ansvarsfördelningen mellan ECB ( Europeiska centralbanken ) , de nationella centralbankerna , kommissionen och Europol ( Europeiska polisbyrån ) vad gäller samtliga frågor som rör förfalskning av euron .
Jag undrar också om det inte vore nödvändigt att upprätta ett interinstitutionellt organ eller EU-organ med ansvar att samordna samarbetet .
Kopplat till detta är också upprättandet av ett system med tidig varning som arbetar dygnet runt , liksom grundandet av ett gemensamt informationssystem för ett snabbt informationsutbyte mellan de ansvariga myndigheterna .
Vid sidan av betänkandet , vilket vi välkomnar , har det dykt upp många frågor som det återstår att reda ut .
Jag hoppas att den diskussion vi för här också skall leda till många klarlägganden .
Herr talman , kära föredragande , kära ledamöter !
Hur säker är euron ?
Detta är en fråga som ju ofta ställs av befolkningen .
Frågan ställs naturligtvis allt mer angeläget ju närmare vi kommer den 1 januari 2002 , det datum då euron kommer att finnas i portmonnän .
Frågan om hur säker euron är gäller nämligen inte endast valutans stabilitet och valutans yttre värde , utan den gäller nämligen även hur man skyddar euron mot förfalskning .
Även detta engagerar befolkningen , för detta penningmedel kommer ju , vilket så riktigt har påpekats , att vara nytt för medborgarna , såväl optiskt sett som när det gäller att handskas med det .
Givetvis blir det även ett nytt faktum för alla medborgare att deras valuta är giltig över ett så mycket större område och dessutom som ledande valuta också utanför Europa .
Även detta är något som man först måste vänja sig vid .
Därför är det klart att frågan ställs vad EU gör för att skydda euron från förfalskning .
Det är också detta det handlar om denna sena timme .
Egentligen är det här en fråga som verkligen står medborgarna nära .
I det hänseendet är det beklagligt att det äger rum så sent på kvällen .
Men det måste ju ske .
Självklart har den Europeiska centralbanken befattat sig med frågan mycket länge .
Centralbanken har ju ansvar för den tekniska säkerheten mot förfalskning .
Kommissionen lade - även det har redan påpekats - sommaren 1998 fram ett meddelande där de mest skilda områden som kräver åtgärder förtecknades , nämligen områdena information , fortbildning - som är en viktig punkt - samarbetet mellan euro-staterna och givetvis samarbetet även utanför detta , samt åtgärderna på straffrättsområdet .
Det är vad föreliggande rambeslut handlar om .
Fru föredragande , jag vill på kommissionens vägnar tacka er så hjärtligt , och framför allt vill jag tacka parlamentet för att ni med så kort varsel var beredda att utarbeta yttrandet .
Det sätter jag verkligen värde på .
I rambeslutet handlar det om att medlemsstaterna skall tillämpa samma definition på valutaförfalskningsbrott .
Det är naturligtvis alltid den första förutsättningen , att man antar samma definitioner för att över huvud taget kunna agera , och det handlar , vilket har poängterats , väsentligen om att skyddet för euron skall garanteras redan innan den existerar fysiskt .
Naturligtvis är kommissionen även tacksam för att Europaparlamentet med sitt snabba beslut - och jag hoppas att det också kommer att röstas så - har gjort det möjligt för rambeslutet att nu träda i kraft så snabbt som möjligt , så att stegen mot ett införlivande nu kan börja tas .
Kommissionen har ju fått i uppdrag och kommer under första halvan av nästa år att lägga fram en rapport om hur det står till med införlivandet i medlemsstaterna , om huruvida allvaret i frågan verkligen återspeglas i motsvarande agerande .
Det har hänvisats till att detta rambeslut är ett beslut på just det straffrättsliga området .
I så måtto måste man godkänna denna reform , denna åtgärd , även om ni , herr Schulz , har påpekat att en komplettering av det tämligen gamla avtalet på det hela taget inte är en alltför djärv åtgärd .
Apropå er fråga om huruvida kommissionen anser att rambeslutet vilar på en tillräckligt stabil rättslig grund i enlighet med fördraget : kommissionen anser att det är rätt grund som tillämpas här .
Emellertid kommer rambeslutet under den närmast följande tiden att behöva kompletteras med ytterligare rättsakter .
Kommissionen kommer att lägga fram ett förslag till förordning om samarbetet mellan samtliga ansvariga myndigheter och om samarbetet med Europol .
Detta förslag skall förpliktiga samarbetet samt reglera de nationella myndigheternas plikt att anmäla fall av valutaförfalskning till Europol samt tillställa Europeiska centralbanken beslagtagna falska pengar för identifikation och klassificering , så att effektiva motåtgärder kan vidtas .
Angående frågan om samordningen av de olika åtgärderna : Sedan början av 1998 arbetar kommissionen och nu i förlängningen OLAF tillsammans med aktuella experter från medlemsstaterna , från Europeiska centralbanken , från Europol , för att på ett effektivt sätt bekämpa förfalskning av euron redan i inledningsskedet .
Från kommissionens sida lades det för några få veckor sedan också fram ett förslag på en informationskampanj om euron - ni , herr Karas , har just påpekat detta - som skall ha en föreslagen finansiering på trots allt 32 miljoner euro .
Detta är ju en finansieringsvolym som kan användas mycket effektivt , dvs. en stor finansieringsvolym ; och givetvis kommer informationskampanjen på en mycket viktig plats även att ta upp eurons säkerhet mot förfalskning .
Och jag tror att den här sena debatten strax före midnatt kan få alla valutaförfalskare på bättre tankar som tror att deras tid är nu , därför att EU inte vakar så sent !
Tack så mycket , kommissionär Schreyer .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
( Sammanträdet avslutades kl .
23.50 . )
