 
Justering av protokollet från föregående sammanträde Protokollet från gårdagens sammanträde har delats ut .
Finns det några synpunkter ?
Fru talman !
Jag vill uttala mig i en fråga som har stor betydelse för alla i denna kammare .
I går eftermiddag svarade kommissionen på frågor under den vanliga frågestunden .
Provan , som var talman , fick stora problem eftersom Byrne använde 29 minuter till att svara på frågor .
Det är särskilt viktigt för denna kammare att vi har möjlighet att ställa frågor till kommissionärerna och jag tycker det är löjeväckande att en kommissionär tar upp 29 minuter för att svara på frågor .
Jag vet att han var särskilt oroad över att behöva svara på en fråga som jag vet att en rad av mina kolleger - inte jag själv - ville ställa till honom rörande skälet till varför han inte vidtog interimistiska åtgärder mot fransmännen i nötköttsfrågan .
Förutom detta vill jag föreslå att - vem som än är talman - om vi får en annan situation då en kommissionär bara pratar på tiden ut , skall talmannen ha befogenhet att stoppa kommissionären eller få honom att korta ned sina svar .
Tack , herr Sturdy .
Jag skall ge ordet till Provan .
Jag vill i förbigående påpeka att han hanterat en något känslig fråga på ett utmärkt sätt , med tanke på hur litet tid vi hade .
Jag tror att för så viktiga meddelanden som detta är en halvtimme verkligen för kort .
Jag tror att vi måste överväga att utöka talartiden .
Fru talman !
Jag är glad att denna fråga tagits upp , men jag hade tänkt ta upp den i parlamentets presidium , vilket är det korrekta förfarandet .
Vi kanske bör ha en diskussion i presidiet om hur vi kan strukturera denna typ av debatt på ett lämpligt sätt i framtiden .
Det var inte tillfredsställande i går .
Vi höll på fem minuter längre än avsett .
Precis som Sturdy sade talade kommissionären i 29 minuter och ledamöterna hade bara sex minuter på sig att ställa frågor .
Det var en löjeväckande situation som vi måste komma till rätta med .
Ja , herr Provan , vi skall granska det vid nästa presidium .
Fru talman !
Ursäkta mig - jag tar sällan till orda i en sådan här situation , men den här gången är det också för att vädja till oss själva .
Trots att jag högaktar Sturdy , uppfattar jag hans klagomål mot Byrne som orättvist ; vi bad nämligen till slut Byrne att presentera vitboken om livsmedelssäkerhet .
Det är en mycket komplex sak som inte kan avhandlas på tio minuter .
Byrne använde 15 till 17 minuter till den , varpå vissa av oss ställde frågor som ibland översteg en minut .
Själv använde jag mindre än en minut , andra mer .
Det är vår uppgift att se till att man inte bara avsätter en halvtimme för kommissionens uttalande , utan en hel timme så att vi har tillräckligt med tid att debattera .
Det Provan sade stämmer .
I går var jag här i plenumet från kl .
15.00 ; det var vi i parlamentet som satte upp oljekatastrofen Erika på föredragningslistan och det var vi i parlamentet som satte upp stormarna i Europa på den .
Allt detta sammantaget ledde till att vi , under vice talmännen Colom och Provan , använt längre tid för våra anföranden .
Det är parlamentet självt som bär skulden för att vi dragit över så pass mycket .
De vice talmännen har inte haft det lätt och det är orättvist att angripa kommissionären för detta , för Byrne fick vänta och blev själv lidande på grund av det .
Det är vi själva som bör ändra föredragningslistan och vara mer disciplinerade .
( Applåder ) Tack , fru Roth-Behrendt .
Ni bekräftar min uppfattning att en sådan debatt egentligen skulle vara berättigad till en dryg timme .
Jag tror att vi kommer att ta hänsyn till detta i framtiden .
Fru talman !
I eftermiddag skall den årliga debatten om inrättandet av området för frihet , säkerhet och rättvisa hållas .
Det är infört i föredragningslistan som frågor till rådet .
Den muntliga frågan skall faktiskt inleda den debatt som förutsetts i utkastet till artikel 2 i fördraget .
Jag vill att ordförandeskapet försäkrar att rådet , som inte har besvarat frågorna skriftligen , i första hand svarar på de frågor som ställts av utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikesfrågor så att vi därefter på ett effektivare sätt kan inleda debatten om EU-fördraget .
Tack , fru Terrón I Cusí .
Vi skall naturligtvis granska detta med rådet .
Vi har gått litet utanför justeringen av protokollet .
Finns det några andra synpunkter på det ?
Fru talman !
Rörande protokoll 21 vill jag att ni noterar vad jag anser vara en tydlig överträdelse av förfarandebestämmelserna i samband med min fråga nr 66 i går kväll .
Den handlar om märkningen av Nestlés bröstmjölksersättningsburkar som tillverkats i Europeiska unionen , vilken skett på ett olämpligt språk och med förvirrande textning och färgsättning , vilket är en tydlig överträdelse av EG : s direktiv 92 / 52 om modersmjölkersättning .
Detta rapporterades först den 5 oktober förra året och såldes fortfarande i Islamabad i Pakistan i går , när jag kontrollerade detta .
Jag vet att ni inte kan kommentera denna fråga rent innehållsmässigt , men genom sitt svar misslyckas kommissionen med att ta ansvar för genomförandet av detta direktiv , på samma sätt som man misslyckats med att tillhandahålla de årliga rapporter som krävs , och som man misslyckats med att följa upp ett tidigare klagomål man fått - se min fråga nr 2283 / 99 .
Jag ber er att skriva till kommissionen på Europaparlamentets vägnar och uppmana denna att fullfölja dess åtaganden , och på vägnar av mödrarna till de 82 barn på varje tusental barn som dör i späd ålder och för vilka användningen av olämplig mat som blandas med orent vatten är livsfarlig .
Helt riktigt , herr Howitt .
Ert inlägg kommer naturligtvis att tas till dagens protokoll , men jag skall också skriva till kommissionen så som ni önskar .
( Protokollet justerades . )
 
Det portugisiska ordförandeskapets verksamhetsprogram samt situationen i Angola Nästa punkt på föredragningslistan är rådets uttalande om det portugisiska ordförandeskapets verksamhetsprogram samt situationen i Angola .
Fru talman , ärade ledamöter !
Det är en stor ära för mig att vara här i Europaparlamentet för att presentera det portugisiska ordförandeskapets verksamhetsprogram för det första halvåret 2000 .
Ledamöterna känner redan till texten i detta program , varför jag kommer att begränsa mig till att betona några av dess viktigaste punkter .
Jag vill börja med att säga att mitt land anser att ordförandeskapets arbete skall bedrivas inte bara med önskvärd effektivitet på ministerrådsnivå , utan också genom ett djupgående samarbete med institutionerna och alla gemenskapsorgan , liksom genom ständig öppenhet i ordförandeskapets verksamhet gentemot den europeiska allmänheten .
Det portugisiska ordförandeskapets förbindelse med Europaparlamentet förtjänar speciell uppmärksamhet eftersom den har en speciell roll inom den interinstitutionella ramen och för att detta organs legitimitet härrör från de europeiska medborgarnas direkta val i de olika länderna .
Detta är det första budskap jag här skulle vilja knyta till löftet om att ordförandeskapet hela tiden kommer att stå till förfogande för klargöranden och ett fullständigt och öppet samarbete med denna kammare .
Fru talman , mina damer och herrar !
Europa befinner sig i dag i ett avgörande ögonblick när det gäller att slå fast den politiska och ekonomiska organisationsmodellen och att fastställa sin identitet på global nivå inför de nya utmaningar som måste besvaras .
Projektet att skapa stabilitets- och utvecklingsvillkor för hela kontinenten , vilket utgör det stora politiska målet för denna europeiska generation , tvingar oss till några val med konsekvenser för unionens framtida projekt .
De senaste åren har vi lyckats uppnå mycket betydelsefulla framsteg när det gäller skapandet av en inre marknad och vi har successivt etablerat det ambitiösa projekt den gemensamma valutan innebär .
Nu måste vi gå ännu längre : vi måste se till att dessa framsteg följs av en parallell utveckling av politiken på andra områden för att ge en fastare struktur åt en enhetlig process som kan svara mot den europeiska befolkningens stora bekymmer och önskningar .
Om vi inte lyckas använda de instrument vi har , det vill säga det Europa som vi har åstadkommit hittills , på ett effektivt och övertygande sätt , är det uppenbart att vi inte kan stimulera våra medborgares vilja att acceptera byggandet av ännu mer Europa .
Det portugisiska ordförandeskapet kommer att försöka se till att den europeiska sociala modellen i framtiden skall utvecklas på ett konkurrenskraftigt sätt och bibehålla unionens förmåga att gå i spetsen för den ekonomiska konkurrenskraften på ett internationellt plan .
I avsikt att stödja förverkligandet av detta projekt , kommer vi nästa månad , i mars , att genomföra ett extra toppmöte med Europeiskt rådet som kommer att ta upp ämnet " sysselsättning , ekonomiska reformer och social sammanhållning för ett Europa med inriktning på innovation och kunskap " .
Det finns säkert några bland er som frågar sig vad vi vill åstadkomma med detta initiativ .
Kan denna tanke tillföra något mervärde till det som redan har gjorts ?
Eller försöker Portugal inleda en ny process som skall läggas till de som utformades i Luxemburg , i Cardiff och i Köln ?
Frågan är befogad och en del av svaret har ni framför er i det dokument som den portugisiske premiärministern offentliggjorde för två dagar sedan .
Det är vår avsikt att med detta arbetsprojekt skapa en bättre förbindelse och samordning av de pågående processerna , genom att även införa en ny dimension .
Vi måste se till att Europa får ett nytt uppsving som gör det möjligt att inom tio år bli det mest dynamiska och aktiva ekonomiska området på världsscenen .
Därför är det viktigt att se till att den europeiska ekonomin lyckas optimera alla sina instrument , och särskilt att den inte släpar efter i den avgörande kampen om konkurrenskraften .
Enligt vår mening går denna kamp via demokratisering av informations- och kunskapssamhället på europeisk nivå , genom att inom detta ämne på ett radikalt sätt minska det avstånd som separerar oss från andra områden som vi konkurrerar med inom den internationella ekonomin .
Denna ansträngning att modernisera , aktualisera och samordna nya resurser avser vi att lägga fram vid Europeiska rådet i Lissabon .
Vi räknar med alla , med detta parlament , med arbetsmarknadens parter , med andra områden inom det civila samhället , och naturligtvis med regeringarna i medlemsstaterna för att kunna genomföra detta viktiga mål .
Fru talman , mina damer och herrar !
Den politiska splittringen på den europeiska kontinenten upphörde redan för några år sedan .
Enandet av Europa har nu blivit det strategiska mål som Europeiska unionen måste arbeta med helt och hållet och som det inte får råda några tvivel om .
Under decennier har det sagts till de befolkningar som har lidit under en begränsad åsiktsfrihet att här , i denna del av Europa , höll en frihets- och framstegsmodell på att skapas som vi önskade att alla skulle kunna delta i .
Nu är tiden inne att visa att vi är konsekventa med det vi har sagt .
Utvidgningsprojektet för Europeiska unionen och alla modeller för avtal som vi avser att skapa med andra länder på kontinenten går i samma riktning : att garantera ett stort område av stabilitet och utveckling som kan ge hela Europa en framtid i fred och framsteg .
Det portugisiska ordförandeskapet har framför sig den viktiga uppgiften att fortsätta de förhandlingar om utvidgningen som inleddes 1998 under stränga tekniska kriterier och en bedömning av objektiva meriter hos var och en av kandidaterna .
Det är vår avsikt att tillsammans med dessa länder öppna alla delar av förhandlingarna i en snabb och effektiv takt , och som grundar sig på förslag som Europeiska kommissionen lagt fram .
Vi kommer på samma sätt att arbeta med fullt engagemang för att ge de sex kandidatländer vi nu börjar förhandla med möjligheten att återta eventuellt förlorad tid utan att detta på minsta sätt påverkar den pågående förhandlingsprocessen .
Det speciella fallet Turkiet kommer att kräva särskild uppmärksamhet från vår sida , med hänsyn till den speciella omständighet som råder och behovet att garantera det land som är en brytningspunkt på världsscenen en fast förhoppning om ett närmande till unionen .
Utvidgningen är alltså ett europeiskt mål som det portugisiska ordförandeskapet inte kommer att undvika utan försöka driva på .
För att utvidgningen skall kunna äga rum anser Europeiska unionen att det är nödvändigt med en reform av institutionerna som gör deras verksamhet mer demokratisk , effektiv och öppen .
Vissa av dessa reformer kan genomföras utan förändringar av fördragen , genom en förbättring av institutionernas arbetsmetoder .
Andra reformer kräver en revidering av fördragen , vilket kommer att ske på den regeringskonferens som vi kommer att presentera inom några veckor , och vi har målet att kunna avsluta den innan detta års utgång .
Det är en erkänt svår och känslig uppgift eftersom den har att göra med beslutsmakten i unionen .
Vår intention är att inviga den med en modell som knyter samman ambition och realism , det vill säga att den lyckas gå så långt som möjligt och nödvändigt med en enhällighet som garanterar att resultaten kan accepteras av medlemsstaterna före slutet av år 2000 .
Respekten för detta är som alla vet , knutet till den omständigheten att varje förlängning av debatten kan leda till förseningar i utvidgningsprocessen , en situation som kommer att få negativa politiska effekter som vi måste ta i beaktande .
Vi är medvetna om att vi med denna nya reform riskerar att inte uppfylla förväntningarna hos vissa och vi känner väl till de befogade önskemål som många i detta parlament har om att gå längre .
Jag kan försäkra att det portugisiska ordförandeskapet kommer att göra allt för att göra agendan för denna konferens , inom det mandat som det fick i Helsingfors , till en samling ärenden som kan utgöra en substantiell reform , men när jag utlovar denna strävan från ordförandeskapet kan jag naturligtvis inte lova några mirakel och speciellt inte att den gemensamma viljan hos medlemsstaternas regeringar skall komma i nivå med era förväntningar och önskningar .
Detta är det sanna och ärliga språk jag här använder inför er , för jag vill inte skapa några falska illusioner .
I detta sammanhang skulle jag vilja ta upp ännu en punkt som oroar det portugisiska ordförandeskapet , eller rättare sagt , som alltid har oroat mitt land , även innan vi övertog ordförandeskapet : Europaparlamentets representation under denna regeringskonferens .
När det gäller denna fråga , som vi också vet är känslig , är vår inställning att , utan att försöka undvika det som är förutsatt i Helsingforsslutsatserna , försöka gå så långt som möjligt med parlamentets deltagande , både i den formella ram som fastställdes i slutsatserna och i de informella modeller där denna institution anser det vara lämpligt med ordförandeskapets samarbete .
Även om vi måste erkänna att vi står inför en representationsmodell som är en förbättring av den status Europaparlamentet hade under förhandlingarna om Amsterdamfördraget , anser vi att det är viktigt att arbeta i en riktning som kan gynna skapandet av en förtroendeingivande stämning och ett effektivt samarbete mellan rådet och parlamentet .
I detta syfte skrev jag till Europaparlamentets talman och meddelade att ordförandeskapet avser att inleda arbetena med regeringskonferensen genom ett speciellt ministermöte vid sidan av rådets ( allmänna frågor ) möte i februari , vilket beslutades i Helsingfors .
Det kommer alltså att bli tillfälle i början av varje ministerkonferens , att utbyta intryck med talmannen och två företrädare för detta parlament .
Detta organ kommer också att ha två observatörer närvarande under alla möten med förberedelsegruppen som kommer att ledas av statssekreteraren för Europafrågor .
Jag tillade i brevet att ordförandeskapet engagerar sig också i att se till att Europaparlamentet får delta på ett effektivt sätt i debatten om regeringskonferensens dagordning .
Vi är öppna för att delta i varje annan arbetsmodell som parlamentet , med respekt för Helsingforsslutsatserna , anser vara lämpligt .
Jag vill försäkra er om att ni kan räkna med oss i detta gemensamma arbete .
Fru talman , ärade ledamöter !
Unionens roll i världen kan bara göra sig gällande i försvaret av dess principer och intressen att göra Europas röst trovärdig , om vi kan åstadkomma ett effektivt svar på de konflikter som uppstår inom strategiska områden och som vi inte kan stå likgiltiga inför .
Kosovokrisen var och fortsätter att vara , möjligen med olika tolkningar , en lektion för oss alla , vilken vi måste dra nödvändiga lärdomar av .
Jag anser att det nu , mer än tidigare , har blivit nödvändigt för Europa att förfoga över egna resurser för att effektivt och i tid kunna agera för att hantera kriser och genomföra operationer för att bevara stabiliteten och freden inom områden som är vitala för vår kollektiva säkerhet .
Europeiska rådet i Helsingfors gav det portugisiska ordförandeskapet i uppgift att genomföra nya säkerhets- och försvarsmekanismer i Europa , förenliga med de åtaganden vissa av oss har inom Atlantpakten , liksom med den speciella situation som drar in vissa partner i Europeiska unionen .
Det är dessutom viktigt att vi kan se till att denna nya modell är helt förenlig med de intressen våra partner i Nato har , både på europeisk och transatlantisk nivå .
Under dessa sex månader kommer vi att pröva den gemensamma viljan att arbeta inom detta område och försöka utforma en enhetlig modell som kan sammanfoga olika ståndpunkter och intressen på ett komfortabelt sätt .
Det är en erkänt besvärlig uppgift , men vi är övertygade om att det handlar om en ytterst viktig utmaning för unionens externa åtgärder , och vi kommer naturligtvis att granska de möjligheter som våra samtidiga ordförandeskap i Europeiska unionen och Västeuropeiska unionen ger oss .
Jag vill också göra några kommentarer om unionens externa förbindelser i mitt anförande , fru talman , ärade ledamöter , och understryka några extra aspekter i det portugisiska ordförandeskapets verksamhetsprogram .
Vi anser att de europeiska ansträngningarna för att få stabila fungerande institutioner inom unionen hela tiden måste ske parallellt med en fortsatt stark uppmärksamhet på det som sker utanför deras område .
Europa har alltid vunnit när det har lyckats underhålla en aktiv och öppen yttre dimension , när det inte flytt in i sig självt för att slippa möta utmaningarna från yttervärlden .
Vi måste nu möta denna värld ansikte mot ansikte och ha en aktiv närvaro i den .
Därför tänker vårt ordförandeskap genomföra en samling åtgärder som främjar och förstärker Europas närvaro i världen , dels genom att följa upp de traditionella förbindelser vi redan har , dels genom att främja nya initiativ inom områden som vi måste sätta i centrum för Europas agenda .
Vi kommer givetvis att rikta särskild uppmärksamhet på den allvarliga situationen på Balkan och på förbindelserna med Ryssland och Ukraina , framför allt på de spänningsområden som påverkar området i närheten av unionen .
Vi strävar också efter att behålla Medelhavsområdet bland våra externa prioriteringar , varför vi kommer att ta flera initiativ i Barcelonaprocessen och försöka få ett synligt engagemang från unionens sida i fredsprocessen i Mellanöstern .
Ett första och viktigt steg togs genom den rundresa jag nyss gjorde i regionen , då jag tillsammans med den höge representanten för den gemensamma utrikes- och säkerhetspolitiken och kommissionen besökte Syrien , Israel , Palestina , Jordanien , Egypten och Libanon .
Det är fortfarande vår intention att utveckla en integrerad politisk dialog med hela Afrika , liksom att garantera att den process som skapats inom området för Lomékonventionen får en tillfredsställande uppföljning i framtiden .
Latinamerika förtjänar en speciell plats inom denna ram för externa åtgärder på grund av den växande betydelse området har för Europa och överensstämmelsen mellan intressen som i dag förenar oss med detta område .
Den transatlantiska dialogen med Förenta staterna och Kanada kommer också att ha en viktig plats på vår dagordning , med hänsyn till det som utgör vårt gemensamma deltagande i de euro-atlantiska institutionerna och särskilt vårt engagemang för att inom den närmaste framtiden , åter få i gång debatten i Världshandelsorganisationen .
Många andra initiativ , framför allt inom en multilateral ram och en bilateral politisk dialog skulle kunna framhävas .
Jag skall dock begränsa mig till att betona den nyhet som toppmötet med Indien kommer att innebära , liksom ministermötena med Australien och Nya Zeeland .
Fru talman , ärade ledamöter !
Jag vill inte dra ut på mitt anförande mer utan lämna tid åt frågor vilka jag med största glädje kommer att besvara .
Jag vill emellertid inte sluta utan att uttrycka två viktiga prioriteringar , som vi kommer att lägga ned arbete på , och en fråga som har direkt samband med arbetet i denna kammare .
Det första spörsmålet gäller det rättsliga området och inrikesområdet : det handlar troligen om en av de expanderande sektorerna i unionens verksamhet som efter Amsterdam har visat sig mer lovande .
På detta område väntar vi på konkreta förslag från Europeiska kommissionen som gör det möjligt för oss att förverkliga ett område med frihet , säkerhet och rättvisa i linje med medborgarnas förväntningar på det europeiska projektet .
Den andra frågan handlar om problemet med livsmedelssäkerhet : vi har just nu en extremt känslig situation på europeisk nivå vilket skapar en stämning av misstroende , med effekter för vår inre marknad , och som på ett negativt sätt projiceras på konsumentskyddet , förutom att det har återverkningar på våra externa förbindelser .
Vi anser att det är viktigt att förändra denna inställning .
Därför är det mycket viktigt att vi lyckas få en enhetlig arbetsram på europeisk nivå , främst genom skapandet av en byrå som kan fungera som ett instrument för samordning av de olika nationella inställningarna .
Det förslag som kommissionen nyligen lade fram , inom ramen för sin vitbok , kommer att behandlas på lämpligt sätt under det portugisiska ordförandeskapet , främst genom en rapport som kommer att läggas fram för rådet i Feira i juni .
Slutligen skulle jag vilja göra klart att frågan om parlamentets ledamotsstadga måste få tillräcklig uppmärksamhet från ordförandeskapet eftersom vi anser det oumbärligt att garantera en viktig aspekt som gäller värdigheten i den verksamhet som utförs inom denna institution .
I detta sammanhang kommer vi att göra vårt bästa för att i dialog med er och i ett gemensamt arbete i rådet , se till att uppnå en rättvis och balanserad lösning på detta problem .
Detta är de viktigaste budskap , fru talman , mina damer och herrar , som jag vill förmedla från den portugisiska regeringen nu när det portugisiska ordförandeskapet för unionen inleds .
Jag står givetvis helt och hållet till ert förfogande för extra klargöranden som ni anser nödvändiga .
Tack så mycket för er uppmärksamhet .
( Ihållande applåder ) Jag tackar rådets ordförande för detta inlägg och jag ger genast ordet till kommissionär Patten , för kommissionens räkning . .
( EN ) Låt mig tacka utrikesminister Gama för hans oerhört tankeväckande och omfattande presentation .
Jag är glad att hans besök i Mellanöstern gick så bra .
Jag är ledsen att jag inte kunde vara där med honom , eftersom jag vid tidpunkten försökte att komma till Thessaloniki för att delta i det första sammanträdet med återuppbyggnadsbyrån .
Jag måste betona ordet " försökte " , eftersom jag under största delen av måndagen befann mig på Münchens flygplats .
Jag har inte för avsikt att tala länge i dag , inte minst därför att jag inte vill förekomma det tal som ordförande Prodi kommer att hålla här nästa månad .
Detta tal kommer inte bara att handla om de kommande sex månaderna , utan de kommande fem åren .
Låt mig emellertid upprepa ordförandeskapets ord och säga att kommissionen naturligtvis kommer att fortsätta att lägga stor vikt vid dess ansvarighet inför detta parlament .
Vi stöder också ordförandeskapets initiativ för att effektivera ministerrådet .
I egenskap av kommission är vi redan engagerade i en omfattande reformering , vilken vi skall diskutera med parlamentet under de närmaste månaderna .
Men jag vill först och främst koncentrera mina kommentarer till frågor som faller under min behörighet som kommissionär med ansvar för yttre förbindelser .
Ordförandeskapet har ett bredare intresse .
Det måste inta en ledande roll under regeringskonferensens första fas .
Det måste också följa upp de många åtaganden som gjordes vid Europeiska rådets toppmöten i Helsingfors och Tammerfors .
Vad gäller t.ex. utvidgningen , kommer formella förhandlingar med de sex nyligen godkända ansökarländerna att inledas i februari .
Samtidigt måste förhandlingsrytmen med de övriga ansökarländerna upprätthållas och föranslutningsstrategin för Turkiet måste upprättas .
Inom alla dessa områden kommer kommissionen att arbeta för fullt .
Andra större initiativ kommer att vara Europeiska rådets toppmöte i mars om sysselsättning , ekonomiska reformer och social sammanhållning för ett kunskapsinriktat och innovativt Europa , och ministern hänvisade till detta .
Vi har för avsikt att följa upp detta toppmöte med en handlingsplan - E-Europa för informationssamhället .
Inom mitt eget område , identifierar ordförandeskapet på ett korrekt sätt utvecklingen rörande formulerandet av den gemensamma säkerhets- och försvarspolitiken som en viktig prioritering .
Minister Gama riktade med rätta uppmärksamheten på betydelsen av att eliminera klyftan mellan Europas ekonomiska styrka och vårt politiska inflytande , inte på grund av någon form av post-imperialistisk högfärd , utan därför att våra medborgare förväntar sig att vi skall göra det och att världen vill att vi skall göra det .
Ordförandeskapet kommer att få se inrättandet av den interimistiska politiska och säkerhetskommittén .
Jag har föreslagit att kommissionen bör skapa ett mindre krishanteringscentrum för att göra det möjligt för oss att reagera snabbare när detta behövs , först och främst rörande biståndsleveranser .
Kommissionen bedömer det också vara viktigt att inrätta en fond som skall utnyttjas när det krävs snabba insatser , och som alltså skall tillhandahålla medel till krisförebyggande åtgärder och krishanteringsverksamhet .
Detta bör t.ex. omfatta ett snabbt utnyttjande av polisstyrkor och mänskliga rättigheter eller övervakare av val , och stöd till civilt biståndsarbete , till säkerhet vid uppbyggande av institutioner och till mediareformer och offentliga informationskampanjer .
Vi kommer även fortsättningsvis att vara engagerade i Balkanområdet och stödja Bernard Kouchner och den FN-ledda förvaltningen i Kosovo , och utveckla våra förbindelser med oppositionen i Serbien för att uppmuntra till ett regeringsskifte , vi kommer också att stödja den demokratiska regeringen i Montenegro , fortsätta den svåra uppgiften med att skapa ett mångkulturellt Bosnien , stödja den nya regeringen i Kroatien och försöka föra Albanien och den f.d. jugoslaviska republiken Makedonien närmare Europeiska unionen .
Låt mig bara ta upp tre allmänna punkter .
För det första måste vi göra allt vi kan för att se till att våra begränsade resurser används på bästa sätt .
Jag har tidigare tagit upp det saktfärdiga och ineffektiva tempot i samband med våra biståndsprogram .
Jag börjar få en stämpel på mig för att vara besatt av denna fråga - en stämpel som jag tycker är hedrande .
Alla som kommer till mitt kontor kan se att mattorna är vältuggade och väggarna välklättrade i frustration över den tid det tar för oss att få saker och ting gjorda .
Det är oacceptabelt - det måste och skall ske en förändring .
( Applåder ) Som jag sagt innan , har jag äran att arbeta med tjänstemän som är mycket bra , men som tvingas följa förfaranden som är usla .
Detta är skälet till varför vi har inlett en granskning av utfallet för våra externa biståndsprogram och jag hoppas kunna lägga fram ändringsförslagen i denna kammare under våren .
Det gläder mig att detta är ett ämne som ni uppenbarligen tillmäter betydelse .
Vi håller på att utarbeta en ny förordning som omfattar vårt bistånd till Balkanområdet .
Avsikten är att förenkla våra förfaranden och påskynda vårt bistånd .
Vi kommer att tillsammans med Javier Solana rapportera till Europeiska rådet i Lissabon om vår politik inom Balkanområdet och bättre sätt på vilka vi kan genomföra vårt bistånd .
I måndags inledde Europeiska återuppbyggnadsbyrån sitt arbete i Thessaloniki .
Den kommer att spela en viktig roll , först och främst i Kosovo och sedermera , förmodar jag , på andra platser .
Jag hoppas den kommer att få möjlighet att följa vår insatsstyrka i Pristina i spåren , vilken nu närmar sig slutet på sitt uppdrag .
Insatsstyrkan har visat att unionen kan utföra ett seriöst , effektivt och snabbt jobb - med rätt ledarskap - med ett minimum av byråkrati och genom att delegera behörighet till personer inom området .
Genom att berömma det arbete som utförts avser jag inte att ge uttryck för tillfredsställelse när det rör situationen i Kosovo .
Det finns enormt mycket för oss att göra där innan vi kan säga att vi uppfyllt våra åtaganden och ideal .
Det finns ytterligare en punkt som är relevant för frågan om resurser .
Medlemsstaterna måste vara beredda att fatta svåra beslut om vad unionen kan och inte kan göra och uppriktigt erkänna att de i bland gör det svårare för kommissionen att vara effektiv , p.g.a. de villkor som lägger sten på börda när det handlar om att genomföra våra initiativ .
Detta kommer att bli ett avgörande år för Ryssland i och med valet av Jeltsins efterträdare .
Tjetjenien kommer naturligtvis att överskugga allt .
Vi kommer ständigt att granska vår politik .
Kommissionen behöver mycket tydliga riktlinjer från medlemsstaterna rörande användningen av de instrument som står till vårt förfogande : Den gemensamma strategin , partnerskaps- och samarbetsavtalet , Tacis , mänskliga rättigheter och demokratiprogram , livsmedelsbistånd osv .
Vi håller på att diskutera med rådet hur vi skall genomföra de beslut som fattades i Helsingfors .
Det kan finnas skäl till att känna sig hoppfull rörande Mellanöstern .
Utvecklingstakten för fredsprocessen i Mellanöstern har påskyndats under den senaste tiden trots bakslag under denna vecka .
Vi kommer inom kort att debattera detta .
Låt mig bara säga att vi är medvetna om att Europeiska unionen måste - vilket också gäller framöver - ge ett större bidrag , och inte bara genom att gräva djupare i våra kollektiva fickor , även om vårt ekonomiska bidrag har varit , och kommer att fortsätta vara , betydande .
I vårt närområde måste vi ge nytt liv åt Barcelonaprocessen , och jag ser fram emot den konferens som kommer att anordnas senare i år om partnerskapet mellan EU och länderna kring Medelhavet , precis som jag ser fram emot toppmötet mellan EU och Afrika .
Jag hoppas att vi skall kunna arbeta med ordförandeskapet vid skapandet av växande politiska och ekonomiska förbindelser mellan Europeiska unionen och Asien .
Kommissionen kommer inom kort att utarbeta ett meddelande tillsammans med Indonesien .
Vi hoppas att våra diskussioner med Kina om inträde i Världshandelsorganisationen ( WTO ) - även om dessa kommer att bli krävande - får att lyckosamt slut .
Det gläder mig mycket att vi , tack vare ordförandeskapets initiativ , kommer att hålla ett toppmöte med Indien .
Jag anser att vi bör arbeta för att stärka våra förbindelser med detta land som ju är den största demokratin i världen ; ett land där - i val efter val - fler röstar i fria och rättvisa val än i hela Europa och Nordamerika tillsammans .
Detta parlament har , förståeligt nog , alltid haft ett starkt intresse av hur Europeiska unionen stöder de mänskliga rättigheterna och demokratiseringen i världen , också genom de hundra miljoner euro som finns tillgängliga inom Europeiska unionens initiativ för demokrati och mänskliga rättigheter .
Jag delar också starkt detta intresse .
Det har skett många förändringar under de senaste åren , inte minst antagandet under 1999 av de två förordningarna med anknytning till de mänskliga rättigheterna .
Under första halvåret innevarande år har kommissionen för avsikt att anta ett meddelande i vilket dess politiska förhållningssätt inom detta område fastställs , inklusive den officiella styrningen av våra program för mänskliga rättigheter och demokratisering .
Parlamentet uppmanade den föregående kommissionen att utvärdera Europeiska unionens deltagande i valobservationsdelegationer under de senaste åren - en erfarenhet som bäst kan beskrivas som " blandad " .
Som svar på denna begäran och på de förändrade rättsliga och budgetmässiga förhållandena enligt de nya förordningarna , har kommissionen för avsikt att anta ett meddelande före påsk , i vilket man kommer att lägga fram vissa förslag till rationalisering och förbättring av vår verksamhet inom områdena valobservation och bistånd .
Jag vet att detta särskilt kommer att engagera denna kammare .
Det kommer helt enkelt att bli mycket jobb de kommande sex månaderna , då vi - hoppas jag - kan få saker och ting gjorda .
Jag ser fram emot att få arbeta tillsammans med kammarens ledamöter och med det nya ordförandeskapet , som jag vill gratulera vad gäller deras program .
Jag ser fram emot att få arbeta tillsammans med dem för att uppnå detta mål .
( Applåder ) Fru talman , herr rådsordförande , kommissionär Patten , kära kolleger !
Såväl rådsordföranden som kommissionär Patten har talat om nödvändigheten av ett gott samarbete mellan institutionerna .
För det vill jag uttrycka mitt eftertryckliga stöd ; jag vill för Europeiska folkpartiets grupps ( kristdemokrater ) och Europademokraters räkning säga att vi eftersträvar ett så nära samarbete som möjligt med rådsordförandeskapet .
Med kommissionen har vi redan ett gott samarbete i allmänhet , och goda kontakter har vi också börjat få .
Det är min förhoppning att vi under det sex månader långa portugisiska rådsordförandeskapet kommer att kunna upprätthålla dessa goda kontakter liksom samarbetet , så att vi i slutändan kan nå gemensamma framgångar .
Framgång för er i rådsordförandeskapet är nämligen också vår framgång - och dessutom framgång för Europa .
Låt oss därför bedriva ett gott och nära samarbete .
Herr rådsordförande , Portugal innehar för andra gången rådsordförandeskapet .
Vi har det största förtroende för er , men se nu till att sätta upp höga mål !
Regeringskonferensen är det största projekt ni kommer att initiera under ert ordförandeskap .
Vi vill bestämt uppmuntra er att prestera ett eget bidrag till fortsättning utöver de tre så kallade leftovers från Amsterdam , och till ett mer ambitiöst program för oss .
Förbered er på att under ert rådsordförandeskap lägga fram sådana förslag som gör att vi kan gå utöver de tre ämnesområdena av leftovers från Amsterdam - toppmötet i Helsingfors ger uttryckligen befogenhet till det , och vi uppmuntrar er till det ; enbart att genomföra dessa tre leftovers är inte tillräckligt för att den kommande regeringskonferensen skall bli en framgång .
Vi måste därför gå längre ; jag vill uppmuntra er att utnyttja er av er rätt att lägga fram nya förslag för regeringskonferensen .
( Applåder ) Jag har nu inte för avsikt att gå in på några detaljer - även om det lockar .
Men sådant hör hemma i debatterna , och mina kolleger Dimitrakopoulos och Leinen har ju lagt fram ett betänkande med en generell inställning som vi delar .
Ställ alltså ambitionerna högt .
Men en sak måste vi självklart se till att hålla hårt på .
På toppmötet i Helsingfors talade man om Europaparlamentets båda observatörer .
Jag ber er av hela mitt hjärta att göra allt som står i er makt under konferensen för att dessa båda företrädare för Europaparlamentet i så stor utsträckning som möjligt får status av likaberättigade deltagare på konferensen , samt även att de förses med teknisk utrustning och arbetsbetingelser sådana att Europaparlamentet kan göra sig hört som anstår det .
Detta vill jag verkligen och av hela mitt hjärta be er om .
Ert rådsordförandeskap lär dessutom faktiskt också bedömas i förhållande till graden av genomförande av denna idé .
Vi vill också tacka kommissionen för att kommissionens ordförande Prodi i Helsingfors gav sitt stöd till vår parlamentsordförande Nicole Fontaines förslag om en bred ansats för regeringskonferensen samt om behovet av att Europaparlamentets båda företrädare får reella möjligheter att delta .
Under det portugisiska rådsordförandeskapet kommer förhandlingar med sex olika länder att återupptas - fem centraleuropeiska länder samt Cypern .
Vi i Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater har alltid begärt att Centraleuropa skall betraktas som en enhet och vi hoppas att man under nästkommande månader kommer att kunna nå framsteg vid förhandlingarna , som lär bli hårda .
Vi ber er också om att ge hög prioritet åt frågorna om den inre säkerheten på den europeiska kontinenten ; dessa frågor är inte bara i sig högst betydande utan de utgör tillika en mycket viktig punkt för acceptansen av utvidgningen i Europeiska unionens medlemsländer .
Ni gav en kort kommentar angående Turkiet .
Europaparlamentet har konstaterat att Turkiet i Helsingfors blivit tillerkänt kandidatstatus .
Vi menar nu att man i den konkreta utformningen av förbindelserna till Turkiet skall tillämpa samma bedömningsgrunder som för de centraleuropeiska länderna .
För att ta ett exempel : Om vi gällande den ungerska minoriteten i Slovakien eller i Rumänien insisterar på att den skall få bevara sin identitet , så förväntar vi oss samma sak från turkisk sida vad gäller hanteringen av kurdfrågan .
På det området vill vi se framsteg så att de etniska minoriteternas identitet kan bevaras även i Turkiet ; vi uppmanar er att vidta motsvarande initiativ .
( Livliga applåder ) Vad gäller Ryssland : Vi behöver stabilitet i Europa .
Vår kontinents säkerhet kommer i stor utsträckning att påverkas av om förhållandena i Ryssland är stabila .
Detta får emellertid inte medföra att vi bara stillatigande åser händelseutvecklingen .
Herr rådsordförande , vi är förpliktade till att göra vår röst hörd med anledning av händelserna i Tjetjenien ; vi måste göra klart för Ryssland att om man fortsätter så här fjärmar man sig från våra europeiska normer om mänsklig värdighet och mänskliga rättigheter .
Var alltså inte alltför diplomatiska när ni tar upp våra betänkligheter mot behandlingen av tjetjenerna och respekten för deras mänskliga rättigheter .
Vi måste göra vår röst hörd .
Kommissionär Patten har med all rätt talat om Medelhavsområdet .
Vår partigrupp är överens om att förbindelserna till Medelhavsområdet , läget i Nordafrika och i Mellersta Östern är lika betydelsefulla för Europeiska unionen som utvecklingen i de centrala och östra delarna av Europa .
Vi tillerkänner det en hög prioritet och eftersträvar en dialog mellan de olika kulturerna .
Men vi vill också be om att man inte har alltför bråttom med att bjuda in vissa personer från Medelhavsområdet till Bryssel .
Man bör nog överväga om inte en sådan inbjudan snarare bör komma mot slutet av fredsprocessen .
Jag skall dock inte fördjupa mig ytterligare i denna fråga .
En avslutande kommentar : Vi har med glädje kunnat höra att ni uttalat er om ledamöternas status .
Parlamentet har lagt fram ett förslag som inte kommer från vår grupp utan från kollegan Rothley , men som vi självklart ställer oss bakom uttryckligen .
Vi vill att en enda rättvis och enhetlig status skall gälla för samtliga ledamöter i Europaparlamentet ; och vi vill värna ledamöternas integritet genom det ; jag välkomnar uttryckligen vad ni sagt om detta - dock måste det vara en enhetlig stadga som gäller för samtliga ledamöter i Europaparlamentet .
Lyckas ni med detta och även övriga programpunkter då är det en stor framgång för Europa och för oss alla - för stabiliteten , säkerheten och demokratin på kontinenten ; vi önskar er lycka till , det här är ingen partipolitisk fråga .
Lycka till från Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokraterna .
( Applåder ) Fru talman , minister Jaime Gama , herr rådsordförande , herr kommissionär , ärade ledamöter !
Jag vill för Europeiska socialdemokratiska partiets grupp hälsa er välkommen , gratulera till ert anförande och till presentationen av det portugisiska ordförandeskapets program och säga att samarbetet med rådet , liksom för övrigt med kommissionen men i detta sammanhang särskilt med rådet , är för vår del inte bara nödvändigt utifrån institutionella kriterier , det handlar om ett samarbete som också krävs i avtalet vi måste respektera på grund av innehållet i det program som det portugisiska ordförandeskapet har lagt fram .
Programmet innehåller en , enligt vår mening , balanserad och ambitiös vision om hur Europeiska unionen bör agera inför de utmaningar vi har framför oss .
Detta sagt om den externa utgångspunkten , med en strategiskt visionär politik i relationerna med flera områden och regioner i världen , och särskild tyngdpunkt på förståelsen av vad som händer i Latinamerika och i Sydamerikanska gemensamma marknaden , men också på prioriteringen av utvidgningen och behovet att fördjupa försvars- och utrikespolitiken i Europeiska unionen .
Men samtidigt som denna vision finns , väl framställd i ordförandeskapets program , finns också en prioritering av och oro inför européernas angelägenheter , inför problem i de länder som utgör Europeiska unionen , med en prioritering av ett område med frihet , säkerhet och rättvisa och även av omsorgen om livsmedelssäkerheten och skyddet för konsumenternas rättigheter och miljöfrågorna , i en vision om hållbar utveckling som bärs upp av detta område självt och inte av någon annan .
Men av alla dessa aspekter , herr minister , är det en sak vi vill ge en eloge för och som är en av det portugisiska ordförandeskapets prioriteringar , det är att man koncentrerar sig på de sociala frågorna och sysselsättningen .
Det portugisiska ordförandeskapet nöjde sig inte med att i sitt program skriva in det som var kvar från andra råd : det valde , det ville göra en markering och en markering som för oss socialister , och säkerligen för majoriteten av ledamöterna i denna kammare , är en viktig markering : inte bara att göra Europeiska unionen till ett dynamiskt och konkurrenskraftigt område på global nivå utan framför allt att vara trogen sina samhälleliga värden och att försvara en europeisk social modell .
Att vara angelägen om en konkurrenskraft grundad på innovation och kunskap är kanske , i början av detta nya årtusende , det bästa bidrag man kan ge Europas grundare och Europeiska unionens verkliga solidaritetsprojekt .
Jag är glad att kunna notera , genom det sätt som dokumentet presenterades på i förra veckan av rådets ordförandeskap och genom dess utformning , att denna punkt kan bli , inte bara en prioritering för ett ordförandeskap , utan också ett signum för Europeiska unionens närmaste framtid .
Vi gratulerar därför till valet av denna prioritering , och vi är beredda att samarbeta för att fördjupa den och för att vi faktiskt skall kunna gå från ord till handling .
Den andra frågan handlar om regeringskonferensen , vilken redan har tagits upp av Poettering .
Europaparlamentet blev djupt besviket på slutsatserna från rådet i Helsingfors .
Besviket på hur rådet ser på Europaparlamentet och besviket på agendan .
När det gäller fördragsreformen vill inte Europaparlamentet förvisas till en roll som observatör av arbetet under denna regeringskonferens .
Vi har åsikter , vi arbetar , vi har erfarenheter och vill bidra med dessa erfarenheter för att hjälpa till så att Europa och Europeiska unionen kan utvecklas och fördjupas ännu mer , och när det gäller dagordningen och dess innehåll , handlar det inte om någon nyck eller halsstarrighet från Europaparlamentet .
Vi tycker inte att man kan ha en regeringskonferens varje år , och vi menar att vi nu har ett tillfälle att föra in några ämnen - inte alla , inte genomföra hela reformen , men föra in några ämnen - , i denna dagordning .
Frågor som försvarspolitiken och medborgarnas rättigheter , vilka kanske behandlas vid sidan om , överenskommelsen om stadgan om grundläggande rättigheter och frågan om en europeisk åklagare är frågor som enligt vår mening , skulle kunna finnas med på denna dagordning , bland andra som kommer att framträda mer i detalj , och därför är jag glad över att notera ordförandeskapets uttalande om att det är för en substantiell dagordningen .
Vi kan kalla den substantiell , global , vi kan ge den fler punkter , men jag gläds åt att notera att det genom seriositet och utan voluntarism , vilket var det uttryck som ministern använde , finns det en beredskap från det portugisiska ordförandeskapet att , tillsammans med Europaparlamentet , kunna få de andra regeringarna att omfatta fler ämnen på denna dagordning .
Detta arbete kan inte bara krävas av det portugisiska ordförandeskapet .
Var och en av oss , i våra länder , var och en av oss tillsammans med kollegerna i de nationella parlamenten har ansvaret för att påverka de andra regeringarna så att vi kan uppnå enhällighet i detta ämne , och den fråga jag skulle vilja ställa , herr minister , är om det kommer att ske några framsteg och om det portugisiska ordförandeskapet , ifall Europaparlamentet kommer med sitt yttrande i tid för att regeringskonferensen skall kunna inledas den 14 februari , redan under det extra Europeiska rådet i Lissabon ämnar lägga fram ett förslag till dagordningen för denna nya regeringskonferens .
Herr rådsordförande !
Jag önskar er lycka till .
Er uppgift är inte lätt , det portugisiska ordförandeskapets program är , som Barón Crespo sade , mycket ambitiöst , men som en gång en portugisisk poet skrev , " när en människa drömmer växer världen och skrider framåt " , och det är när det finns höga ambitioner som man kan ta steg framåt , även om det skulle vara små steg , mot att göra Europeiska unionen starkare , mer solidarisk och framför allt mer förankrad hos alla dess medborgare .
( Applåder ) Fru talman , herr rådsordförande , herr kommissionär !
Jag vill ta tillfället i akt och på ELDR-gruppens vägnar lägga fram tre förslag till det tillträdande ordförandeskapet .
Låt mig först säga vad gäller utvidgningen , att vi verkligen välkomnar förändringen i vad som jag skulle beskriva som " stämningen " och de politiska ambitionerna kring utvidgningsdebatten .
Detta bekräftades i Helsingfors och det ligger nu i ordförandeskapets händer att utveckla detta material .
Rörande de ansökarländer som redan börjat förhandla är det tydligt att vi nu börjar närma oss de mer kritiska och komplicerade delarna av förhandlingsprocessen , och för de som just fått klarsignal i Helsingfors måste vi nu inleda detta arbete med .
I detta sammanhang är det viktigt att uppmärksamma och ta itu med vissa av de element som tydligt håller på att växa fram inom den allmänna debatten .
Det är tydligt att det i vissa ansökarländer finns en viss avmattning hos allmänheten rörande det europeiska projektet .
Det är viktigt att uppmärksammar och tar itu med detta i det politiska arbetet .
I vissa fall finns det tecken på en framväxande " de och vi " mentalitet , och vi måste ta itu med denna .
Jag vill föreslå ordförandeskapet att ni förutom de vanliga diplomatiska kanalerna , genom vilka ni i ert uttalande om mål åtagit er att rådfråga ansökarländerna om deras planer och regeringskonferensen , bör överväga att använda den europeiska konferensen som en mekanism och en metod att på ett offentligt sätt lyssna och delta i en dialog med ansökarländerna om deras synsätt .
Vi föreslår detta som ett medel att på högsta politiska nivå demonstrera den likhet som råder rörande bedömningen av ansökarländerna .
Min grupp anser att det är viktigt att man engagerar sig i att skapa ett partnerskap för Europa och inte ett Europa som skapas genom diktat .
Vi måste hitta mekanismer för att tydligt få våra ansökarländer att förstå detta under förfarandets gång .
Den andra fråga som jag vill ta upp handlar om regeringskonferensen .
Det åvilar er att genomföra den oerhört viktiga uppgiften att fastställa dagordningen och starta konferensen - i bland tror jag att det är en ganska otacksam och svår uppgift .
Det är tydligt att konferensen kommer att handla om det som blev kvar efter toppmötet i Amsterdam .
Detta är naturligtvis viktigt , men jag menar att det inte är tillräckligt vad gäller en ambitiös inställning till dagordningen och jag delar de åsikter som andra kolleger som talat i dag har framfört .
Man kan nästan känna det kyliga draget av den stängda dörren i Helsingfors om frågan rörande mer långtgående ambitioner , men slutsatserna lämnade emellertid denna dörr på glänt .
Herr rådsordförande !
Jag vill uppmana er att på ett bestämt sätt placera er fot i dörrspringan och förespråka en mer ambitiös dagordning .
Det är oerhört viktigt att vi nu tar tillfället i akt genom denna regeringskonferens och försöker att ge tillbaka litet själ till Europa .
Det är mycket tydligt att fördragens nuvarande konstruktion misslyckas med att på ett meningsfullt och tillgängligt sätt fånga strävandena i vårt samtida Europa .
Fördragen misslyckas med att på ett tydligt och heltäckande sätt visa för en vanlig person hur institutionerna fungerar .
Vi måste bli bättre på att förklara detta genom att bygga in det i de grundläggande dokumentens struktur , och jag ber er att börja om från början .
Det kanske var för tidigt att utropa ett ambitiöst " ja " i Helsingfors .
I dag är det för tidigt att säga " nej " .
Börja om från början med detta , så får ni denna kammares stöd .
Jag välkomnar verkligen ert engagemang i samband med denna idé om ett innovativt och kunskapsinriktat Europa och jag ser fram emot att bidra till denna debatt i denna kammare och direkt med ordförandeskapet .
Vi har utfört mycket arbete tillsammans med Förenta staterna om den digitala dialogen , för tillfället i synnerhet inom områdena rörande privatliv och dataöverföring , men det är inte slutfört .
Vi har ett lagstiftningsforum mellan denna kammare och den amerikanska kongressen .
Vi har regelbundna toppmöten mellan rådet och Förenta staterna och det finns allt färre möjligheter att avsluta vissa fall med en avgående förvaltning .
Jag uppmanar er , herr rådsordförande , att ta kontroll över denna dagordning och dra vissa specifika och tidiga slutsatser av den transatlantiska digitala dialogen och inte låta den flyta bort för att återupptas på nytt vid ett senare datum av en annan förvaltning .
Det är nu den verkliga möjligheten finns och ni kan slussa igenom den som en del av ert initiativ rörande ett innovativt Europa .
Kör hårt och lycka till !
( Applåder ) Herr rådsordförande !
Genom en lycklig omständighet i tidsplanen får ni ta över ett särskilt ansvar : inleda en regeringskonferens som uppenbarligen är grundläggande för Europas framtid .
Ni kommer också - och det är den andra frågan jag skall ta upp - att vara ordförande för en konferens vars betydelse inte undgår någon , om sysselsättning och ekonomisk och social sammanhållning .
När det gäller regeringskonferensen vill jag gärna berätta om min grupps ståndpunkt och även om vilka förslag vi har .
Innehållet till att börja med - olika kolleger som talat har med rätta betonat att Helsingforsmötet var otillräckligt , och en så snäv föredragningslista förefaller oss inte godtagbar .
Vi vill absolut att minst fyra konkreta punkter skall tas upp på dagordningen : juridisk status för stadgan med de grundläggande rättigheterna och dess inverkan på medborgarna , det förstärkta samarbetet som är en grundläggande mekanism , den successiva integrationen av utrikes- och säkerhetspolitiken , med särskild betoning på förebyggande av konflikter inom gemenskapspelaren och slutligen översyn av det ålderdomliga Euratomfördraget , som bör ses över när det gäller målsättningarna och sedan införlivas i unionens fördrag .
När det gäller metoden har regeringskonferensens åtgärder länge tydligt visat sina begränsningar , liksom regeln om enhällighet .
Rådet gjorde misstaget att inte ändra metod .
Vi är besvikna över det men om rådet vill visa att man vill ha en mer demokratisk och starkare union , måste man åtminstone ta med Europaparlamentet så mycket som möjligt , och jag vill också lägga till de nationella parlamenten .
Europaparlamentet bör på samma sätt som kommissionen vara delaktigt , eftersom vi är de två institutioner som har en gemenskapsvision , och det skulle vara logiskt att parlamentet blir delaktigt i ett samtyckesförfarande i slutet av förhandlingarna .
Annars är jag , liksom andra kolleger , rädd att gapet vidgas mellan allmänheten och de europeiska institutionerna .
Vi upplevde i Seattle ett viktigt förfarande , en livlig reaktion från det civila samhället gentemot en världsomspännande institution som man inte förstår och vars funktion uppfattas som farlig för samhället i sin helhet .
Det får inte bli på samma sätt för Europeiska unionen , det skulle jag personligen beklaga .
Ni skall snart resa runt i huvudstäderna för att övertyga era kolleger om att man skall utvidga dagordningen och ändra metoden .
Vi avvaktar resultatet av era åtgärder innan vi uttalar oss om framtiden för denna regeringskonferens .
Jag skulle slutligen vilja betona en punkt som enligt min uppfattning inte förts fram tillräckligt : det är i stort sett nödvändigt att lyckas med konferensen annars riskerar vi att definitivt blockera Europeiska unionen .
Jag tänker på ett område som ligger oss varmt om hjärtat , nämligen skattefrågan .
Sedan flera år är vi inte i stånd att fatta ambitiösa beslut om skatter på miljöområdet , eftersom enhällighetsregeln hindrar oss från det , och jag kommer nu till den andra punkten i mitt inlägg , nämligen sysselsättningen , eftersom denna typ av beskattning också kan generera sysselsättning .
När det gäller toppmötet om sysselsättningen har man talat om innovation och alla är positiva till det .
Även om innovation definitivt kan öka konkurrenskraften , får man ändå inte skyla över en verklighet som är mindre lysande och mer oroande .
Förvisso är det ofta så att innovationen spelar en viktig roll , men konkurrenskraften förvärvas ibland genom tvivelaktiga mekanismer : en i vissa fall omfattande försämring av arbetsvillkoren i Europa , ökade risker , försämrad miljö och allmän stress .
Det är inga uttalanden tagna ur luften : en rapport nyligen från Europeiska fonden för förbättring av levnads- och arbetsvillkor i Dublin visar att arbetsvillkoren är dåliga eller försämras för ett stort antal arbetstagare ; när det gäller miljön visar 1999 års rapport från Europeiska miljöbyrån att av 12 studerade parametrar motsvarar 11 antingen status quo eller en försämring .
Oljefartyget Erikas förlisning visar för övrigt att konkurrenskraften inom en ekonomisk sektor kan uppnås till priset av försämrade arbetsförhållanden , ökade risker och ett allvarligt hot mot miljön .
Jag tror därför att det är på tiden att se över vissa gällande mönster och jag beklagar att det inte framgår tydligare av ert dokument .
Jag tror exempelvis att innovation kan kombineras med en strävan efter att öka inte arbetets produktivitet utan produktiviteten av sällsynta resurser och icke förnybara resurser .
Det är säkert en utmärkt väg att gå , inte bara för en hållbar utveckling utan också för att skapa sysselsättning som är stabilare , säkrare , mindre stressande och mer lovande för framtiden .
Vi kommer nu tillbaka till utgångsläget i mitt inlägg .
Allt detta kan bara ske om vi förändrar de europeiska institutionerna .
Det är därför den målsättning vi måste satsa på .
Fru talman , herr rådsordförande !
Jag vill välkomna det portugisiska ordförandeskapet och säga att vi mycket uppmärksamt kommer att följa de vägar som tas angående detta ordförandeskaps viktigaste frågor och prioriteringar : från utvidgningen till fördragsrevisionen , från Lomékonventionens framtid till toppmötet Europa-Afrika , från sysselsättningsproblemen till de som gäller andra och tredje pelaren .
Vi kommer att göra detta främst på grund av de farhågor som några av dem väcker , eller kanske det sätt de tas upp på .
Detta är fallet med utvidgningen , vars förverkligande vi inte har några principiella skäl emot , men vars genomförande vi anser oansvarigt , om det sker utan en djupgående analys i förväg av olika konsekvenser och hur man skall förekomma dem .
Till detta kan nu läggas ännu större farhågor inför att Turkiet räknas som kandidatland , när vi fortfarande bevittnar dess regerings totala ovilja att lösa kurdfrågan på ett adekvat sätt eller att upphöra med ockupationen av Cypern .
Även revideringen av fördragen väcker allvarliga farhågor .
Inte så mycket på grund av en möjlig och effektiv anpassning av dessa till utvidgningen , utan för att vi befarar att man , med detta som förevändning , skall falla för frestelsen , och det oacceptabla misstaget , att skapa en politisk ledning för Europeiska unionen .
När det gäller Afrika tar vi med en blandning av tillfredsställelse och viss oro emot meddelandet , som inte bekräftades av ordförandeskapet här , om att dörrarna åter står öppna för genomförandet av det toppmöte som sedan tidigare har planerats .
Tillfredsställelse eftersom vi alltid ansett det nödvändigt och lägligt att förverkliga det , särskilt om det inriktas på ett verkligt samarbete mellan de två kontinenterna , enligt lämpliga modeller , men också för att vi alltid har hävdat att vi måste fortsätta att göra allt för att kunna genomföra det .
Dock även med en viss oro eftersom det presenteras med mycket kort framförhållning , till april månad , som är den planerade tidpunkten för toppmötet , vilket säkerligen gör det svårt att planera mötet på lämpligt sätt , om det inte till och med äventyrar dess genomförande .
Vi noterar därför på vederbörligt sätt ordförandeskapets nya uttalande om Angola .
Trots att det är sent från rådets sida , tycker vi att det går i rätt riktning , även om vi , framför allt i ljuset av de ståndpunkter vi själva har intagit här i parlamentet och i den gemensamma församlingen , hade hoppats på en mer fördömande inställning av UNITA med tanke på dess otvetydiga ansvar för hela det drama landet upplever .
Men lika mycket som , eller mer än , formen för vissa frågor som står i fokus under det närmaste halvåret , oroas vi av det faktum att vissa frågor som är avgörande för oss , inte finns med bland det portugisiska ordförandeskapets prioriteringar .
Den ekonomiska och sociala sammanhållningen glöms bort , och anses nästan diabolisk på gemenskapsnivå , och det är tråkigt att behöva konstatera att även det portugisiska ordförandeskapet undviker att alls nämna främjandet av sammanhållningen , trots att ordförandeskapet innehas av ett av länderna med lägst relativ utveckling .
Det låga valdeltagandet i de senaste valen till Europaparlamentet bekräftade det djupa demokratiska underskottet och visade på medborgarnas stora avstånd till de dominerande nyliberala inriktningarna .
Trots detta , och trots att vi står inför en fördragsändring , ser vi inte några institutionella förändringar som kan göra slut på detta underskott , och under tiden insisterar man på dessa inriktningar utan att göra något för att framför allt bekämpa arbetslösheten på ett effektivt sätt och främja sysselsättningen , frågor som är mycket angelägna för medborgarna .
Genomförandet av ett extra toppmöte om ett pompöst ämne lugnar oss inte , eftersom vi redan har haft flera toppmöten om sysselsättningsproblemen utan att det lett till någon vilja att förändra den dominerande penningpolitiken , och även därför att målen och tidsfristerna är så vaga och ambitionerna med programmen motsägelsefullt oproportionerliga och tycks snarare vara en rökridå än en händelse med verkliga avsikter att förändra gemenskapens status quo på ett påtagligt sätt .
Herr rådsordförande !
Vi kan i dag analysera det program som har lagts fram och avsikter med detta .
Men i juli kan vi göra en noggrann fullständig slutbedömning av det portugisiska ordförandeskapet , och det kommer vi att göra .
Fru talman , herr minister och rådsordförande , herr kommissionär , kära kolleger !
Det roterande ordförandeskapet är ett av de mest unika kännetecknen för Europeiska unionen .
Varje halvår är det som om vi alla står inför en ny inledning och återigen drar oss till minnes den eviga andan , samma eviga anda , varken mer eller mindre .
De inriktningar som har fört oss hit , som har åstadkommit det som hade varit otänkbart för femtio år sedan , är samma grundläggande inriktningar - dessa och inte andra som vi har velat skapa - som dessa och andra framtida förenta stater i Europa kan föra ännu längre .
Det är klart att känslan av att börja om mycket är en illusion .
Kontinuiteten i våra ärenden kan inte ta någon hänsyn till olika Europa var sjätte månad , men det är en mekanism som friskar upp minnet genom nya infallsvinklar och påminner oss om vad vi är : ett Europa med partnerskap mellan länder , ett nationernas Europa .
Jag hoppas att förväntningarna på det portugisiska ordförandeskapet uppfylls vad gäller ett kreativt och varaktigt sammanfogande av arbetena i Luxemburg , Cardiff och Köln , och i förbindelserna med Afrika , och i arbetet med moderniteten - informationssamhälle och digital-TV - eller i omsorgen om gemenskapens yttersta randområden .
Jag tror att vi i allmänhet borde vara djärvare i befästandet av framtiden för den ekonomiska och sociala sammanhållningen , ett centralt mål för fördragen , långt ifrån uppfyllt , vilket också är bland dem som mest attraherar utvidgningsländerna .
När regeringskonferensen sätter i gång rekommenderar vi försiktighet och realism .
Den fråga som debatteras i Europa i dag är deltagandet : ett effektivt deltagande från befolkningarna , i linje med de verkliga känslorna hos allmänheten i länderna .
Det låga valdeltagandet i valen till Europaparlamentet har diskuterats flera gånger .
Det är ett problem som inte påverkar parlamentets legitimitet , men som pockar på en demokratisk ödmjukhet från oss alla , och får oss att avstå från en våldsam förvandling av unionens karaktär eller fördragens struktur och balans .
Mer än att förvandla allt , bör vi förbättra det vi har , och börja här i denna kammare , i vårt sätt att debattera , genomföra omröstningar , hur vi förmedlar det , hur vi kommunicerar och umgås med våra kolleger i de nationella parlamenten , och det är också rekommendabelt med en viss blygsamhet .
Därför håller jag inte med om muttrandet om att parlamentets yttrande skulle fördröjas i reaktion mot en åberopad brist på stadga .
Detta vore en allvarlig ansvarslöshet och det är inte problemet .
Problemet , för det handlar om fördragsrevideringen , är det bristande deltagandet från de nationella parlamenten innan , ett område där vi med intresse kommer att följa inriktningen på ordförandeskapets program .
Problemet här är att det bara finns en observatör från de två största politiska grupperna i stället för en från varje konstituerad grupp .
Problemet med deltagande löses genom att utvidga deltagandet , inte genom att insistera på ännu fler av samma Dupont och Dupont .
Jag vill inte sluta utan två oumbärliga anmärkningar om två färska händelser .
Jag vill inte i dag , som portugis till portugis , kalla det kritik , snarare en nödvändig oenighet .
För det första , en oenighet med beslutet att inte förlänga vapenembargot mot Indonesien .
Det är ett olyckligt beslut och mycket olägligt .
Det verkar som om vi glömmer bort de döda som fortfarande håller på att begravas i Östtimor , den osäkerhet som fortfarande består och det cyniska dubbelspel de indonesiska militära myndigheterna spelar .
Det som vi alltid har kritiserat har skett : en total svaghet i ett beslut som har fattats på sikt i stället för med tydliga villkor .
För det andra , en oenighet också vad gäller uttalandet om Angola .
Det är ytterliga en olycklig händelse .
Det är ofullständigt , obalanserat och hjälper inte fram någon lösning på en långvarig tragisk konflikt .
Vi stöder inte heller UNITA : s agerande de senaste åren , men det innebär inte att ansluta sig till krigets väg , att strunta i de mycket allvarliga anklagelserna om en fruktansvärd krigsekonomi som skadar den angolanska staten , att ta ställning för ena parten , att assistera eller till och med samarbeta i plundringen av resurser till olycka för en befolkning som är drabbat av ett krig sedan decennier , att ge kritikerna rätt i att utländska aktörer agerar på ett oacceptabelt partiskt sätt .
När det gäller Angola kan målet bara vara ett : fred , medlen kan bara vara ett fåtal : fredliga och dess uttryck kan bara vara ett : en humanitär radikalism .
När det gäller det lidande som drabbar befolkningen har ingen av de krigförande parterna i Angola rätt .
Det har de inte !
I vilket fall som helst , efter denna nödvändiga parentes önskar jag det portugisiska ordförandeskapet all framgång .
Herr Gama !
Vi gläds åt ert ordförandeskap som inleder årtusendet , eftersom ni i Bryssel med de aktuella och brådskande frågorna om Timor och Macao , meddelade oss vad som kunde bli Europas öde : att ha varit och inte längre vara .
Tidsplanen ger er av en tillfällighet en roll som ni känner till väl , eftersom er namne Vasco da Gama också var upptäckare .
Ni skall öppna vägen mot regeringskonferensen .
Men först har vi de återstående ärendena , såsom samarbetsavtalet med Sydafrika och det särskilda avtalet om vin : porto , ouzo , grappa och sherry piratkopieras av Sydafrika och Sydafrika kommer inte att respektera sitt åtagande .
Vad tänker ni göra ?
Bland de andra återstående ärendena har vi också euron ; euron fungerar som gemensam valuta .
Varför ändra en situation som fungerar ?
För mervärdesskatten har övergångsperioden behållits .
Varför inte göra samma sak när det gäller euron ?
Utöver det stora antalet ärenden har vi det sociala toppmötet om sysselsättningen i mars .
Om inte ett mirakel sker som i Fatima , om man inte ger sig på den överdrivna internationaliseringen och de överdrivna skatterna , kommer man inte att lösa problemet .
Vad tänker ni göra åt det ?
Sedan har vi regeringskonferensen .
Vi avvaktar med ångest dess resultat , särskilt som vissa vill inrätta en europeisk åklagare .
Ni kommer att göra rättvisan till en prioriterad fråga .
Ni har hos er Sid Ahmed Rezala , mördaren som Frankrike släppt ut , som Spanien befriat och som nu är hos er .
Vi får väl se vad ni beslutar att göra med honom .
Slutligen har vi öppningen mot öst , i väster börjar Europa hos er .
Hur långt går det i öster ?
Fram till gränsen mot Iran , till Kaukasien , från Lissabon till Moskva ?
Herr Gama !
Ställ de rätta frågorna på alla dessa punkter .
Vi får väl se om era franska socialistkamrater som efterträder er lämnar de rätta svaren .
Fru talman !
Det finns nu en tidtabell för mer union , men det vi har behov av är en tidtabell för mer demokrati .
Den 10 februari kommer Portugal att lägga fram ett förslag till dagordning för regeringskonferensen .
Den 14 februari inleds konferensen .
Den 24 februari sammanträder utrikesministrarna , och därefter sammanträder de varje månad för att diskutera åtminstone fem viktiga frågor .
För det första har vi frågan om majoritetsbeslut .
På hur många av de 65 områden som vi i dag har ett förfarande med enhällighetsbeslut kommer det framöver att vara majoritetsbeslut , så att demokratierna i våra medlemsstater kan röstas ned av ministrar och tjänstemän bakom stängda dörrar i Bryssel ?
För det andra har vi kommissionens sammansättning .
Det kommer nog även framöver att vara en kommissionär för varje land , men de små länderna kommer oftast att få en junior-portfölj .
För det tredje har vi röstviktningen i ministerrådet , parlamentets sammansättning och domstolen .
De fem största länderna får kanske 25 procent fler röster i rådet , även om alla förlorar lika mycket genom utvidgningen .
För det fjärde kommer det att ske ett förstärkt samarbete .
Portugal och andra federalistiska länder kommer att pressa på för att en majoritet av medlemsstaterna skall kunna bygga ut samarbetet , även om vissa länder skulle vara emot , och i detta förhållande ligger det ett faktiskt avskaffande av vetorätten i viktiga frågor .
För det femte finns det en restavdelning som kommer att handla om allt det som medlemsstaterna skickar in , och på toppmötet i Porto kommer man alltså att kunna utvidga dagordningen för det som beslutades på toppmötet i Helsingfors .
Allt kommer att sluta med ett nytt unionsfördrag som skall ersätta Amsterdamfördraget före år 2003 .
Det kommer att antas i Nice den 8 december i år , med det blir knappast nice , om inte väljarna blandar korten på nytt .
Det uppmanar vi gärna till från Gruppen för demokratiernas och mångfaldens Europa , som är min grupp här i parlamentet , och från vår gemensamma tvärpolitiska grupp med meningsfränder som heter SOS Demokrati , för det är SOS Demokrati vi behöver , inte mer byråkratmakt i Bryssel .
Herr talman !
Jag vill börja med att tacka rådsordföranden för hans principförklaringar , framför allt beträffande Europaparlamentets medverkan .
Utan tvivel har han en svår uppgift och frukterna av sitt arbete kommer han själv knappast att kunna skörda - det tycks vara ordförandeskapets eviga väsen .
Om jag nu håller mig enbart till problemet med regeringskonferensen så visar enbart diskussionen om föredragningslistans omfång på de stora meningsskiljaktigheter som råder mellan medlemsstaterna .
Med risken att upprepa mig och med vetskap om att jag därmed befinner mig i konflikt med merparten av ledamöterna i kammaren , insisterar jag på att rådets anspråkslöshet i Helsingfors var riktig .
Alla har vi när allt kommer omkring tvingats uppleva hur man i Amsterdam sköt upp och lämnade de frågor som skulle vara regeringskonferensens kärnfrågor utan lösning .
Europaparlamentets katalog av önskemål berör tveklöst flera viktiga frågor .
Dessa önskemål bör emellertid inte tas upp förrän olika leftovers fått sin lösning i stället för att öppna för möjligheten att de viktigaste frågorna återigen förbigås i förhandlingarna .
Först när man lyckats knäcka dessa nötter finns möjligheten att ägna sig åt övriga frågor .
De visionärer som sätter tempot före grundligheten gör mig bekymrad .
Herr talman , minister Jaime Gama , rådsordförande som jag hjärtligt välkomnar , kommissionärer , ärade ledamöter !
I det roterande ordförandeskapet har turen detta halvår kommit till Portugal .
Detta system garanterar en jämlikhet i varje medlemsstats bidrag till det europeiska bygget , om ordförandeskapet genomförs på ett effektivt sätt och att man försöker finna en klok balans mellan nationella krav och uppfattningen av Europas allmänna intressen .
Det är uppenbart att rotationen gör att de viktigaste delarna av arbetet sker enhälligt mellan medlemsstaterna och medborgarna i dessa .
Om inte detta sker , får vi en rad ordförandeskap som inte förstår varandra och som saknar riktlinjer eller styrs av en osynlig hand vilket är oacceptabelt .
Jag hoppas mycket av det portugisiska ordförandeskapet .
Jag hoppas att det skall hjälpa till att svara på den centrala politiska frågan : vart går Europeiska unionen och på vilka vägar ?
Bara då kan vi gå över till den institutionella reformen , vilket är ett villkor för eller en konsekvens av utvidgningen som måste ske i respekt för balansen mellan Europeiska unionens nationer , befogenheter och politik vilken mödosamt har följts under årtionden .
Att bygga upp är svårt och mödosamt , att förstöra går snabbt , vilket motiverar en stor försiktighet i behandlingen av denna fråga .
I denna fråga kan en upplösningsprocess av Europeiska unionen börja .
Några kanske tänker : detta är komplext och väldigt ambitiöst , varför Portugal ?
Jag svarar : om det måste genomföras , varför inte Portugal ?
När det viktigaste är beslutat blir det en del av övriga ärenden .
Det vi anser om Europeiska unionen är oförenligt med vissa lösningar .
Jag kan inte acceptera att man talar om utvidgning till varje pris , så som vissa , kanske för många , gör .
Jag kan inte acceptera att man i en omfördelning av makten , och frågan är huvudsakligen den om makten , överlämnar den till en styrelse som utgörs av de starkaste länderna eller att bara dessa skall få plats och makt i Europeiska kommissionen .
Jag kan inte acceptera att mitt språk inte skulle vara officiellt språk .
Jag kan inte acceptera ett nedmonterande av den gemensamma jordbrukspolitiken eller att den skall fortsätta att gynna några och glömma andra , liksom jag avvisar att solidariteten bryts i sökandet efter en reell konvergens av utvecklingsnivåerna .
Den ekonomiska och sociala sammanhållningen , en fördragsprincip , måste återigen finnas med i första ledet av unionens angelägenheter och prägla alla politikområden .
Jag kan inte acceptera bevarandet av det nuvarande finansieringssystemet , liksom jag inte kan acceptera avsaknaden av en gemensam utrikes- och säkerhetspolitik .
Det talas mycket om medborgarnas Europa .
Man vill ha deras medverkan och informera dem , mobilisera dem kring starka idéer , motsvara förväntningar om genomförande .
Det är inte med en status som mindre värd , vilken Europeiska rådet ger Europaparlamentet under regeringskonferensen , som man erkänner dess representativitet .
Liksom man inte genom att en månad besluta tvärtemot vad Europaparlamentet ansåg månaden innan , kommer att nå framgång : detta inträffade i frågan om vapenembargot mot Indonesien .
Men hur skall man väcka intresse hos medborgarna som många gånger vänder ryggen till ?
Låt oss försöka ge ett svar .
Tillsammans med mina landsmedborgare , ser jag på Europeiska unionen från dess västra gräns i Azorerna , en av de regioner som i Fördraget om Europeiska unionen betecknas som " yttersta randområden " .
Det jag därifrån vill se är lika möjligheter , tillnärmande av de livsvillkor som fortfarande finns där .
Jag ser inte utvidgningen som bara en addering av områden för att motsvara externa politiska utmaningar , jag vill se fördelning , solidaritet , samma förmåga till självförverkligande där jag bor , i norr , öst , syd som i mitten .
Liksom jag är intresserad av de stora frågorna och anser att fördragen har ett perspektiv där människor räknas , följer jag uppmärksamt effekterna av Europeiska unionens små beslut angående min region , som är stor , alltså för mina medborgare .
I detta ögonblick vill vi veta vilka åtgärder man planerar för gemenskapens yttersta randområden .
Vad är framtiden för den mjölkproduktion som vår ekonomi är beroende av , en produktion som sker under unika villkor och som vi vet hur vi skall framställa i en nästan perfekt symbios med naturen ?
Som ni ser hoppas jag mycket av det portugisiska ordförandeskapet .
Jag hoppas att det hjälper till att staka ut en väg och bibehålla den känsliga balansen , och att man i detta sammanhang gör framsteg i mycket viktiga frågor och med egna kännetecken .
Jag hoppas att man engagerar medborgarna , och uppmärksammar deras legitima önskemål .
Jag hoppas att ett arbete för Portugal är ett arbete för Europeiska unionen .
Herr talman !
En av de största utmaningarna som det portugisiska ordförandeskapet står inför är regeringskonferensen .
Som ni känner till mycket väl är detta parlament missnöjt med den tänkta dagordningens inskränkthet .
De tre s.k.
" Amsterdamresterna " är mycket viktiga och omfattar vad som förmodligen är den enskilt mest viktiga frågan för regeringskonferensen i samband med utvidgningen , dvs. den ökande volymen beslut som skall fattas genom ett förfarande med kvalificerad majoritet .
Det är visserligen sant , men dessa tre frågor är mycket välkända för våra medlemsstater .
De har ingående granskat dem under förhandlingarna i Amsterdam .
De känner exakt till frågorna .
De behöver inte granska dessa under ett helt år .
De behöver en överenskommelse .
De behöver förhandla en natt , kanske en vecka , och ett paket att avtala om .
Då återstår resten av året - nästan ett helt år .
Det är dubbelt så lång tid i jämförelse med den regeringskonferens då man ingick avtal om Europeiska enhetsakten 1985 .
Det är lika lång tid som den regeringskonferens då man ingick avtal om det mycket omfattande Maastrichtfördraget .
Denna regeringskonferens varade ett år .
Det är därför fullt möjligt att ta upp andra frågor .
Ingen vill egentligen ha en allomfattande regeringskonferens med hundratals frågor - med en julgran där alla hänger upp sina favoritdekorationer .
Det vi ber om är helt enkelt att ett begränsat antal viktiga frågor skall tillfogas dagordningen ; frågor som man faktiskt borde ta itu med under det som är den sista regeringskonferensen före utvidgningen - sista gången vi har dessa förhandlingar utan att det blir nästan 30 medlemsstater kring bordet , vilket gör alla avtal mer komplicerade än vad som är fallet just nu .
Vi måste ta tillfället i akt .
Det skulle vara höjden av oansvarighet att inte göra det .
Under toppmötet i Helsingfors fick ni - det portugisiska ordförandeskapet - ett mandat att föreslå ämnen som kan tillfogas dagordningen .
Detta innebär , med Cox ord , att dörren står på glänt - liberalerna stjäl alltid de bästa uttrycken från andras tal .
Vi har för avsikt att på ett bestämt sätt placera vår fot i dörrspringan och se till att den fortsätter att stå på glänt och t.o.m. öppnas ännu mer .
Gudskelov för att dörren står på glänt , därför annars hade detta parlament nästan med säkerhet frestats att yttra sig negativt om regeringskonferensens sammankallande , eller t.o.m. att fördröja vårt yttrande och därigenom fördröja starten på regeringskonferensen ; kanske t.o.m. att återkalla våra företrädare från regeringskonferensen .
Men det faktum att dörren står på glänt innebär att det fortfarande finns en väg framåt .
Det som förändrar saken enligt min grupp , är den attityd som uppvisats av det portugisiska ordförandeskapet .
Ni delar tydligen vår oro över dagordningens inskränkthet .
Ni skulle tydligen också föredra att dagordningen utvidgades och ni har gett oss ett löfte att ni skall göra ert bästa i detta avseende , precis som ni just nu har sagt till oss att ni skall säkerställa vidast möjliga tolkning av åtagandena från Helsingfors rörande parlamentets deltagande i regeringskonferensen .
Detta förändrar verkligen saken , vad min grupp anbelangar .
Vi välkomnar detta .
Men just som min kollega , Seguro , vill jag be er att tydligt uppge att ni har för avsikt att lägga fram förslag till en utvidgning av dagordningen redan till Europeiska rådets första sammanträde i Lissabon i mars , och inte vänta till juni .
Detta skulle vara mycket viktigt för att hjälpa till med att övertyga detta parlament att avge sitt yttrande i tid , så att ni hinner inleda regeringskonferensen på alla hjärtans dag den 14 februari .
Herr talman , herr rådsordförande och herr kommissionär !
Det portugisiska ordförandeskapet har onekligen en hel del att göra under våren , inte minst vad gäller arbetet med regeringskonferensen och utvidgningen .
Det kan inte ha undgått er att detta parlament vill se en utvidgad agenda med avsevärda institutionella reformer till fromma för ett mer effektivt och demokratiskt EU .
Om detta kan man tala länge och mycket .
Jag vill dock ta upp en annan fråga som av outgrundlig anledning hamnat på denna punkt på föredragningslistan .
Jag vet att den är angelägen för Portugal , och den oroar min grupp , den liberala gruppen , mycket .
Vi ser med förfäran på den förvärrade situationen i Angola .
Med stigande oro har vi sett hur UNITA-gerillan ökar sina militära aktiviteter och urskillningslöst ger sig på civila , nu senast genom massakern på över hundra civila i Bieprovinsen .
Vi ser också med stor oro på hur yttrandefriheten i landet stryps .
Minst tjugo journalister arresterades förra året , trots att regimen i Angola försäkrat att den respekterar pressfriheten .
Det finns flera enskilda journalister som på minst sagt tvivelaktiga grunder väntar på rättegång , anklagade för förtal av presidenten .
Vi hoppas att de kan få en öppen , rättvis och snar rättegång .
Folket i Angola har alltför länge plågats av detta tröstlösa inbördeskrig som har orsakat tusentals döda , lemlästade , undernärda och över två miljoner hemlösa .
Situationen för civilbefolkningen är akut .
EU har ett historiskt engagemang i Angola och är en stor biståndsgivare .
Det är hög tid att tillsammans med FN öka pressen på Savimbi att återuppta de havererade fredssamtalen , men också pressen på regimen att den måste sluta med sina plundrarfasoner och respektera yttrandefrihet och mänskliga rättigheter .
Vi liberaler utgår från att dessa frågor kommer att ha hög prioritet i samband med Portugals arbete med det nya partnerskapet mellan EU och Afrika .
Herr rådsordförande , herr kommissionär , herr talman !
Ett litet land är vant vid att ha mycket utland och det är lovande , bland annat för de frågor som togs upp av den föregående talaren .
Det sätt på vilket er befolkning , herr rådordförande , har engagerat sig i Östtimor , väcker hoppet att ni skall kunna lägga en grund för ny fred och nytt samarbete i Afrika .
Vi var verkligen besvikna över Helsingfors och den begränsade dagordningen för regeringskonferensen och vi hoppas att ni skall utvidga den maximalt och använda den till förmån för ett starkare samarbete .
I dag och i framtiden måste Europa kunna fungera som en demokrati .
Det går inte utan reformer .
Då blir en utvidgning det samma som en urvattning av unionen .
För vår grupps räkning och särskilt för Europeiska fria alliansen vill jag be om ert ordförandeskaps uppmärksamhet för de regioner och kulturgemenskaper som visserligen inte är medlemsstater men som har grundlagsenlig behörighet för vissa ärenden som de måste kunna samarbeta med Europa om .
Herr rådsordförande !
Vi yrkar för att det skall kunna ske direkt .
Till vår besvikelse togs det i Helsingfors , ett land som ändå är känt för att förorda insyn och öppenhet , ett steg i motsatt riktning i den ökända bilaga 3 .
Jag vill också peka på att vi den här veckan i parlamentet talat om de stora skillnaderna i välfärd mellan regionerna i Europa .
Arbetslösheten i våra fattigare regioner blir knappast mindre .
Hur skall vi kunna förverkliga utvidgningens stora ambitioner om vi inte ens i Europa självt kan uppbringa någon respekt för kulturer , för språk och inte ens kan minska de stora skillnaderna i välfärd mellan våra regioner ?
Jag vet att ni anser att det här är mycket viktigt och jag önskar er stor framgång med det .
Herr talman , herr rådsordförande !
Jag skulle först av allt vilja lyckönska er till ett initiativ från det portugisiska ordförandeskapet .
På ett relativt signifikativt sätt har ingen kollega talat om det , det gäller det första toppmötet Europa-Indien .
Jag anser att det är ett grundläggande initiativ .
Kollegerna föredrar , som de gjorde med Sovjetunionen , att fortsätta att i dag diskutera med Kina , som för övrigt flertalet västföretag håller på att dra sig ur .
Vi fortsätter att främja den röda mattans politik och fjäska för Peking , och vi ser inte att vi kan skapa ett strategiskt avtal med Indien såsom ni vill göra .
När det gäller regeringskonferensen tycker jag att Poettering visade prov på humor i förmiddags när han sade att om de tre leftovers kunde lösas under det kommande rådet blir det en framgång för Europeiska unionen .
Man måste verkligen vara närsynt för att inte inse att om vi inte tar oss an den grundläggande frågan , den om det konstitutionella medbeslutandet , om vi inte kan tänka oss en mekanism som är värdig en parlamentarisk dialektik , kommer vi att med 28 , 30 eller 32 medlemmar snabbt bli fullständigt förlamade .
Jag vill därför uppmana er , herr rådsordförande , att inte alltför noggrant notera denna mycket långa lista med så många punkter som ett stort antal kolleger skulle vilja lägga till en annan lista , som ni för övrigt redan känner till , utan om möjligt begränsa er till att föra in denna enda punkt som kan garantera att Europeiska unionen inte blir förlamad i morgon .
Till de kolleger som förväntar sig ett svar från er när det gäller de två lobbyister som vi redan har vid regeringskonferensen tror jag att det också där är på tiden att vi inser att det inte är med lobbyister som vi kan förstärka en institutionell dialektik , utan att det är vår skyldighet att kräva att Europeiska unionen grundas på verkliga parlamentariska mekanismer , med en dialektik mellan detta parlament och rådet som är värdig namnet , och inte längre små segrar som ger mer eller mindre marginella poäng på regeringskonferensens föredragningslista .
Herr talman !
Portugal har som första ordförandeland för EU det här årtusendet ställt upp ett klart och tydligt verksamhetsprogram .
Ändå har jag några frågor som jag gärna skulle vilja få klarhet i från ordförandeskapet .
För det första är jag glad över att Portugal fäster stor vikt vid den kommande utvidgningen av Europeiska unionen .
Det ger också utrymme till utvidgning av dagordningen för nästa regeringskonferens .
Förutom de tre leftovers från Amsterdam så behövs långtgående reformer för att kunna välkomna de nya medlemsstaterna .
Dessutom prioriterar ordförandeskapet en förstärkning av GUSP .
Förra veckan visade det sig i det gemensamma mötet med den amerikanska kongressen och Europaparlamentet att man även från amerikanskt håll oroar sig över finansieringen av GUSP .
Kommer den att ske på bekostnad av den budget som EU-länderna nu ger till Nato ?
Ordförandeskapet föreslår ett extra toppmöte om bland annat sysselsättningspolitiken .
Jag upprepar vår synpunkt att den mycket hellre kan utformas på lokal nivå .
När det gäller de ekonomiska reformerna så vill jag ta upp Irland och Nederländerna som exempel .
Dessa länder har nu fått ordning på det hela och förtjänar att få efterföljare .
Angående livsmedelssäkerhet står det en hel del i verksamhetsprogrammet .
Men precis vad är det egentligen som ordförandeskapet vill ?
Slutligen undrar jag hur ordförandeskapet hoppas uppnå enighet om stadgan och hur det ser på den oberoende expertundersökning angående tyngden av EP-medlemskap .
Kommer ordförandeskapet att försvara undersökningsresultaten i rådet ? )
Herr talman , herr rådsordförande !
Regeringskonferensens dagordning är inte tillräcklig .
Kommissionen har sagt det och de politiska grupperna i parlamentet har sagt det .
Den är otillräcklig , men slutsatserna från Helsingfors lämnar vägen öppen för en ändring .
Det portugisiska ordförandeskapets uppgift är enligt min mening att försöka åstadkomma en sådan ändring , vilket jag uppmanar ordförandeskapet att göra .
Uppgiften är inte överambitiös .
Det är en uppgift som grundar sig på sunt förnuft .
Vi vill att regeringskonferensen även skall ta upp andra frågor just därför att vi inte vill ha regeringskonferenser vart tredje eller fjärde år .
Vi vill att den här regeringskonferensen skall lösa frågorna för en lång tid framöver .
Herr talman , vi menar att det i huvudsak är tre frågor som borde ingå i regeringskonferensens agenda .
Den första har att göra med Europas roll i världen .
De institutionella aspekterna av säkerhets- och försvarspolitiken , som man under senare tid har gjort stora framsteg med och som en majoritet av européerna stöder , är en fråga som till slut måste tas upp i Nice .
En annan fråga som vi måste reflektera över är det förstärkta samarbetet .
Utvidgningen , vårt mål för de nästkommande åren , Europeiska unionens historiska utmaning , kommer att kräva flexibla formler vid genomförandet av vår politik .
Rättfärdigandet tror jag vi alla känner till .
För att underlätta utvidgningen måste vi därför beakta det förstärkta samarbetet i dagordningen .
Avslutningsvis kan jag nämna en annan fråga som jag också anser vara viktig .
För ett par veckor sedan inledde vi något som i de europeiska medborgarnas ögon är av särskilt stor vikt .
Europeiska unionens dokument om de grundläggande rättigheterna .
I Tammerforsslutsatserna nämns möjligheten av ett uttalande eller att man skall ta med det i fördraget .
Jag tror att vi till slut kommer att vara tvungna att inkludera dokumentet om de grundläggande rättigheterna i fördraget .
Gör vi det uppnår vi något viktigt : en förening mellan Europeiska unionen och medborgarna .
Jag säger det på ert vackra språk genom att citera en portugisisk poet - förena de mänskliga rättigheterna med det där " comboio de corda que se chama o coração " ( " pulserande tåget som kallas för hjärta " ) .
Herr rådsordförande , ni har viktiga uppgifter att ta itu med och parlamentet litar på att ni klarar av det .
Seguro , vår kollega från Europeiska socialdemokratiska partiets grupp , ställde en öppen fråga till er och även jag skulle vilja höra det portugisiska ordförandeskapets svar på denna .
Herr talman , herr rådsordförande , kära kolleger !
Det portugisiska ordförandeskapet har lagt fram ett ambitiöst program .
De europeiska socialisterna litar på Antonio Guterres och hans medarbetare när det gäller att återföra vår union på vägen mot en hållbar ekonomisk utveckling .
Europa lider av flera stora brister .
Vi har fortfarande för hög arbetslöshet .
Vi har en lägre andel sysselsatta än Förenta staterna och Japan .
I Europa är de offentliga och privata investeringarna otillräckliga .
Den nödvändiga budgetkonsolideringen har fått många stater att minska sina investeringar i infrastruktur , men den privata sektorn har inte alltid tagit över .
De s.k. " riskkapitalinvesteringarna " är dubbelt så stora i Förenta staterna som i Europa .
Amerikanerna investerar tre gånger mer än européerna i skapandet av nya företag .
I Förenta staterna går 80 procent av riskkapitalet till ny teknik , jämfört med bara 27 procent i Europa .
Japan investerar 2,9 procent av sin BNI i forskning och utveckling , Förenta staterna 2,8 procent och Europa bara 1,8 procent .
Forskarna utgör bara 2,5 procent av arbetskraften i våra företag , mot 6 procent i Japan och 6,7 procent i Förenta staterna .
Vi lider brist på hjärnor .
Vi har färre universitetsstuderande än amerikanerna och japanerna .
Nära hälften av de europeiska studenter som doktorerar i Förenta staterna stannar kvar där och arbetar .
På teknikområdet finns det 700 000 till 800 000 lediga jobb i Europa , i brist på kvalificerad personal .
Amerikanerna har samma problem .
Förra året inrättade emellertid den amerikanska senaten en kvot på nära 500 000 immigrationsviseringar på fyra år för s.k. högt kvalificerade arbetstagare .
Europa kan inte arrangera en sådan brain drain , en sådan stöld av hjärnor .
Vi måste i stället investera i information , utbildning och innovation .
Innovation och kunnande är i dag de viktigaste källorna till rikedom för nationerna .
Vi måste lyckönska det portugisiska ordförandeskapet till att kämpa för ett Europa av innovation och kunnande .
Rådets ordförande har just aviserat att det inte blir någon Lissabonprocess .
Det är lovvärt .
Vi måste i stället samla processerna från Luxemburg , Cardiff och Köln i en enda samordnad åtgärd med precisa och kontrollerbara målsättningar .
Tillväxt- och stabilitetspakten från Dublin är mycket stabil men innehåller ingen tillväxt .
Stabiliteten är nödvändig , men är inte ett mål i sig och när världens ekonomiska framtidsutsikter ser bättre ut , kan vi hoppas på en Lissabonpakt för sysselsättningen från det portugisiska ordförandeskapet .
Herr talman !
Jag vill här visa min uppskattning för att det portugisiska ordförandeskapet med en sådan handlingskraft tar tag i förberedelserna för den kommande regeringskonferensen .
Det är verkligen goda nyheter efter de inte särskilt tillfredsställande resultaten av toppmötet i Helsingfors .
Min grupp anser att dagordningen för regeringskonferensen måste utvidgas så att Europeiska unionen verkligen skall kunna fungera effektivt med över 20 medlemsstater i framtiden .
Därför är vi glada över att ordförandeskapet vill inrätta fem arbetsgrupper som skall undersöka de viktigaste problempunkterna .
Men liksom många har betonat så är de tre leftovers från Amsterdam en alldeles för mager dagordning .
Min grupp kräver också att Europaparlamentet skall vara en fullvärdig part vid förhandlingsprocessen , vilket Fontaine och andra tidigare med eftertryck har begärt .
Under de kommande veckorna kommer ordförandeskapet att besöka alla huvudstäder i våra EU-medlemsstater .
Vi kräver att det portugisiska ordförandeskapet vid den rundresan till alla huvudstäder i de olika medlemsstaterna i EU utvidgar regeringskonferensens dagordning i enlighet med rekommendationen i betänkandet av Dimitrakopoulos-Leinen .
Jag anser att det portugisiska ordförandeskapet efter den rundresan skall rapportera om resultatet av dessa samtal under sammanträdesperioden i Strasbourg i februari .
Jag skulle vilja påminna ordförandeskapet om att det i artikel 48 i Fördraget om Europeiska unionen står att regeringskonferensen inte kan inledas förrän Europaparlamentet yttrat sig .
Jag utesluter inte att Europaparlamentet ger sitt yttrande först efter att det står klart hur Europaparlamentet på ett bättre sätt skall engageras i förhandlingarna och dagordningen har utvidgats .
Herr talman !
Det ämne som kommer att tas upp i mars är av mycket stor betydelse .
Vi får dock inte inskränka det till demokratiseringen av informationssamhället .
Låt oss främst se efter var Amerika är bättre än Europeiska unionen och inom det området lära oss best practices av Förenta staterna .
Herr talman !
Jag skulle vilja fokusera på sysselsättning och sociala frågor .
Jag välkomnar verkligen det dokument som utarbetats av ordförandeskapet denna vecka , som en del av förberedelserna för det särskilda toppmötet i mars .
Det visar ett berömvärt , sammanhållet förhållningssätt , ett övergripande förhållningssätt som är mycket välkommet - än mer därför att det tar hänsyn till en rad av de viktiga förslag som vi har lagt fram i denna kammare under de senaste åren .
Dessa omfattar behovet av att förbättra samordningen mellan sysselsättningsstrategin och de breda ekonomiska riktlinjerna .
Jag ser fram emot genomförandet av de förslag ni kommer att anta i mars och hoppas att ni får det stöd ni behöver .
Endast en sak gjorde att min glädje inte blev fullständig och det var i samband med konvergensen av social trygghet .
Många av oss i denna kammare hoppades att få se ett Luxemburgliknande förfarande om konvergens av social trygghet , men jag är rädd att texten i dokumentet inte är i närheten av detta , utan i stället talar man om gemensam analys , samarbete och utbyte av bästa metoder .
Detta är inte är inte tillräckligt för att skapa den modernisering av de sociala trygghetssystemen som vi behöver i Europeiska unionen .
Om jag får ta upp specifika sociala paket , finns det två stycken jag kort vill nämna något om .
Ett som är mycket viktigt för oss är de allmänna ramarna om information och rådfrågning .
Jag hoppas att det kommer att ske framsteg rörande detta paket under det portugisiska ordförandeskapet .
Men vi har också moderniseringen av företagsrådsdirektivet , dess granskning och ändringar .
Under de senaste månaderna har jag fått besök av arbetare från Michelin i Frankrike , Ford i Portugal , i går av arbetare från ABB-Alsthom som påverkats av sammanslagningen , arbetare som förvägrats sina rättigheter enligt företagsrådsdirektivet .
Detta måste moderniseras och genomföras av kommissionen .
Kommissionen misslyckas med att uppfylla sina åtaganden .
Om vi är seriösa när det gäller partnerskap på arbetsplatsen och de förbättringar som detta kan medföra ; om vi är seriösa när det gäller innovation och produktivitet , måste vi granska lagstiftningen inom detta område och se till att industrins båda sidor visar lämplig respekt för varandra under denna partnerskapsprocess .
Herr talman !
Herr rådsordförande , ni har lagt fram flera mycket ambitiösa projekt .
Min grupp skulle gärna se att ni också kunde genomföra en stor del av dessa , särskilt på den inre säkerhetens område .
Jag vill framhålla två punkter vilka förefaller mig vara speciellt betydelsefulla .
För det första : Optimeringen av Schengensystemet , säkrandet av de yttre gränserna .
För det andra : Förbättrad asylpolitik samt kampen mot laglöshet och människohandel .
Till att börja med tänkte jag berätta om en aktuell situation i Belgien och vid de belgiska yttre gränserna .
Situationen är bekant : I Belgien infördes helt plötsligt över en natt kontroller av landets inre gränser , vilket medförde timslånga köer och även problem i gräns- , person- och godstrafiken ; detta innebar förtret för medborgarna och störningar på ekonomin .
Skälet var den förestående legaliseringen av ca 75 000 illegala invandrare , som fortfarande , efter tre-fyra års vistelse i Belgien , väntar på besked i asylfrågan eller som redan har fem-sex år av olaglig vistelse i landet bakom sig .
Det kan vara värt att påpeka att åtgärderna som Belgien vidtagit är i enlighet med lagar och fördrag .
Härav blir det dock uppenbart att detta inte kan vara lösningen på de återstående problemen , utan att vi här måste söka oss nya vägar och att lösningen till syvende och sist bara kan göras på gemenskapsnivå .
För övrigt har Belgien valt en väg som liknar den som tidigare Frankrike , Italien och Luxemburg valt .
Ansvaret ligger hos rådet .
Det är anledningen till de krav vi kommer med .
Vad jag vill och vad vi vill är att ni optimerar Schengensamarbetet som ett instrument för säkerheten , att ni företar en förnyad reglering av kontrollerna av de inre gränserna vilka tillfälligt återinförts samt att medlemsstaterna får information på förhand , varvid också tidsutdräkten bör anges ; dock bör detta endast göras i absoluta undantagssituationer ; då måste det dessutom genomföras snabbt och fullständigt över hela gemenskapen .
Det andra är naturligtvis införandet av enhetliga och snabba asylförfaranden , varvid ett omgående införande av Eurodac ter sig som särskilt brådskande ; detta innebär att medlemsstaternas ansvar slås fast och att verksamma instrument mot olagligheter ställs till förfogande .
Herr talman , mina ärade damer och herrar !
Nu skulle jag förstås helst ta upp de förväntningar på rådsordförandeskapet som min kollega Pirker redogjort för .
Det vore roligt , men tyvärr är ju tiden för den typen av diskussioner rätt begränsad i det här parlamentet .
Jag måste av den anledningen skjuta på det till i eftermiddag .
Då skall vi nämligen tala om årsrapporten för området säkerhet , frihet och rättvisa .
Jag vänder mig till det portugisiska rådsordförandeskapet med följande begäran : Det var rådet - inte rådsordförandeskapet - som vägrade att ge parlamentet en skriftlig rapport för utvärdering av utbyggnaden av området säkerhet , frihet och rättvisa .
Det finns en muntlig fråga , dock inget skriftligt svar från rådet ; det motiv man ger till detta är att det inte är tillräckligt om rådet framför detta svar här i dag muntligen .
Förfaringssättet är typiskt inte för rådsordförandeskapet utan för tjänstemännen i rådet , vilka förhåller sig till parlamentet som en överhetsstat .
Överhetsstaten tenderar att säga : Vi , företrädarna för överhetsstaten , bestämmer vad som är bra för folkrepresentationen och vad som inte är det .
Detta har vi i parlamentet ofta fått uppleva inom området säkerhet , frihet och rättvisa .
När vi i morse fick höra det portugisiska rådsordförandeskapets ord att man är beredd att just på nämnda område inleda ett konstruktivt samarbete med Europaparlamentet , så kan vi bara säga att vi verkligen välkomnar det .
Överhuvudtaget menar jag att allt som framförts av det portugisiska rådsordförandeskapet visar på en stor öppenhet gentemot den parlamentariska instansen i Europeiska unionen .
Och det är bra , för vi måste ha klart för oss - speciellt när det gäller den mellanstatliga handeln , som fortfarande finns med i fördraget och fortfarande gäller vid uppbyggnaden av området säkerhet , frihet och rättvisa - att Europaparlamentet kommer att spela en central roll just på de områden där den mellanstatliga handeln äger rum och har omedelbara konsekvenser för de enskilda medborgarna samt mindre medverkan från de nationella parlamenten än tidigare .
Om nu rådsordförandeskapet påstår att man erkänner detta - så har vi förstått det från det portugisiska rådsordförandeskapet - anser jag att vi i parlamentet kan inte annat än ge vårt stöd till det och säga : Om bara alla rådsordförandeskap agerade så , vore kontakterna mellan parlament och råd fungera betydligt bättre på den här nivån .
Herr talman !
Jag vill börja med att välkomna rådets tjänstgörande ordförande och ställa tre betydelsefulla frågor om de utskott i detta parlament som jag sitter med i .
Den första frågan handlar om beslutsprocessen inom den gemensamma jordbrukspolitiken , vilken bara ger Europaparlamentet en marginell funktion som simpel rådgivare .
Vid en tidpunkt då den gemensamma jordbrukspolitiken alltmer betraktas som landsbygdspolitik , den första pelaren i det europeiska området , skyddet av miljön , arvet och sysselsättningen , är det obegripligt att parlamentet fortfarande bara har en rådgivande roll , vilket dessutom innebär att man inte har beslutsbefogenheter för mer än 40 procent av unionens budget .
Den andra frågan handlar om behovet att skynda på genomförandet av den nyligen meddelade europeiska myndigheten för livsmedelssäkerhet .
Men det är viktigt att klargöra om vi bara bryr oss om den europeiska organismen för utvärdering och förvaltning av riskerna eller om vi bryr oss om en substantiell förstärkning av den gemensamma kvalitets- och säkerhetspolitiken för livsmedel , inklusive veterinärernas verksamhet .
Om det är så måste medlen påtagligt ökas , såväl på unionsnivå som på nationell nivå .
Om nu det senaste alternativet gäller , vilket jag anser bör vara fallet , måste jag säga att jag inte lugnas av Europeiska kommissionens meddelande förra veckan , där synen tycks vara att skapa " ytterligare " ett vetenskapligt organ helt utan befogenheter och isolerat från en gemensam åtgärd på alla fronter och länkar i jordbruks- och livsmedelskedjan .
Den tredje frågan jag skulle vilja ta upp handlar om fiskeavtalet mellan Europeiska unionen och Marocko .
Jag oroas verkligen över kommissionens sena inledning av förhandlingarna , liksom över den långsamhet vi kan bevittna från rådets sida i processens framskridande .
Jag måste också säga att jag oroas över att inte i någon del av det portugisiska ordförandeskapets program ha sett ett påskyndande av förhandlingarna om avtalet nämnas .
I gengäld har jag i samma program sett ett omnämnande av att fördjupa analyserna av kostnads- och intäktsanalyserna beträffande fiskeavtalen med tredje land vilket är det argumentet som vanligtvis åberopas i Europeiska unionen av dem som motsätter sig fiskeavtalen mellan unionen och tredje land .
Jag skulle därför vilja höra vad ordförandeskapet har att säga om de frågor jag nu har ställt .
Herr talman , herr rådsordförande , kommissionär Patten , mina damer och herrar !
Jag har det senaste portugisiska ordförandeskapet från 1992 i gott minne .
Under det antogs normer och jag önskar er , herr ordförande , liksom oss alla att ert ordförandeskap blir lika framgångsrikt den här gången .
Ni har lagt fram ett omfattande och ambitiöst program .
Jag skulle vilja sätta fingret på en utrikespolitisk och en säkerhetspolitisk aspekt av programmet och ställa några frågor i anslutning till dem .
Får jag be er att ge detaljerade svar på dessa frågor .
För det första : Turkiet .
Jag har ända sedan början stött Turkiets kandidatur och gläder mig nu över resultatet från mötet i Helsingfors .
Kommer nu ordförandeskapet att stödja denna kandidatur genom att formulera en åtgärdskatalog och en tidsplan och därigenom göra det möjligt för Turkiet att på samma sätt som övriga tolv kandidater komma till förhandlingsbordet ?
Och är ordförandeskapet villigt att ta initiativ för att lösa kurdproblemet ; kanske kan man ge sitt stöd till en konferens på samma sätt som skedde i Madrid för Mellersta Österns vidkommande - här avser jag den idé som Poettering , som tidigare tagit upp kurdproblemet , lanserade ?
Beträffande den gemensamma säkerhetspolitiken ger toppmötena i Köln och Helsingfors anledning till hoppfullhet .
Nu måste något konkret göras .
Det måste vara något som accepteras av samtliga EU : s medlemsländer och som kan accepteras även av de länder som inte är medlemmar i Nato .
Jag har , herr rådsordförande , känslan att ni orienterar er mot Nato och frågar er hur en konstruktion som passar in i Nato kan se ut .
Men det handlar inte om det .
Vad vi behöver är en europeisk konstruktion , som passar ihop också med Nato - det måste vi se till .
Herr talman !
Det portugisiska rådsordförandeskapet har en svår uppgift att tampas med .
De båda föregående rådsordförandeskapen har formulerat mål och slagit fast mandat som kanske inte är särskilt långtgående .
Er uppgift är nu att genomföra detta .
Det kan hända att resultatet i slutändan blir lyckat , men hur som helst är det ni fått på er lott ingen lätt uppgift .
Det gäller särskilt den sista punkten som kollegan Sakellariou tog upp , nämligen frågan om förverkligandet av en europeisk utrikes- och säkerhetspolitik .
Europaparlamentet kommer härvidlag att ge sitt oinskränkta stöd till er ; vi lägger naturligtvis också vikt vid att funktionen som komplement till Nato behålls samtidigt som européerna utvecklar en egen kapacitet på det här området för att därigenom kunna hantera de svåra situationer som kan uppstå .
Ni har också i fortsättningen uppgiften att tillse att Barcelonaprocessen fortskrider ; vidare innebär utvecklingen av förhandlingarna i Mellersta Östern helt nya chanser .
Jag har fått intrycket att de berörda parterna i dag i mycket större utsträckning än tidigare är villiga att acceptera att Europa spelar en roll på detta område .
Jag önskar er och Patten all framgång med denna uppgift .
Ytterligare punkter av vikt är naturligtvis regeringskonferensen , spänningsförhållandet mellan utvidgning och handlingsförmåga i Europeiska unionen samt de problem som kan uppstå i samband med riskerna för overstretching och de nödvändiga beslut som vi måste träffa på regeringskonferensen .
Ni är bunden till ett visst mandat .
Å andra sidan visar erfarenheten att , när en av de parter som deltar i förhandlingarna väl presenterat ett förslag , är det mycket svårt att stoppa en diskussion om förslaget .
Detta innebär att såväl hittillsvarande praxis som era faktiska handlingsmöjligheter ger er möjligheten att tolka mandaten mycket vitt .
Jag tror att förutsättningarna för att vi i Europaparlamentet skall kunna fatta rätt beslut i vårt yttrande är goda , om ni kan ta initiativ till en sådan bred tolkning av mandatet .
Därigenom skulle det i högre grad bli möjligt för oss att lägga fram våra föreställningar om demokrati och Europeiska unionens handlingsförmåga på förhandlingsbordet .
Herr talman !
Efter att ha hört så många ambitiösa och betydelsefulla saker sägas om utrikespolitik och sysselsättningspolitik skäms jag nästan att komma med klagomål .
Men jag måste ändå göra det .
Jag har läst ert verksamhetsprogram och lyssnat uppmärksamt på er .
Jag skulle önska att programmet var lika ambitiöst på de områden jag arbetar för här i parlamentet , nämligen områdena miljöpolitik , konsumentskydd och hälsopolitik .
Jag är medveten om att ett ordförandeskap inte kan ta sig an allt och inte satsa på alla områden , och därför respekterar jag att ni fokuserar på annat .
Men jag kan ändå inte låta er slippa undan så lätt - det förstår ni nog också .
Jag vill göra några kommentarer .
I ert skriftliga program - och även i det som ni framfört här i dag - har ni lagt vikt vid livsmedelssäkerheten .
Det är viktigt .
Parlamentet kommer att ta itu med vitboken " Livsmedelssäkerhet " .
Ministern har påpekat att toppmötet i juni skall befatta sig med den vitboken .
Jag hoppas att ni har så pass stor respekt för Europaparlamentet att ni inväntar parlamentets samråd och även besluten , men jag betvivlar att så blir fallet ända fram till juni .
Vi vill dock gärna göra ett försök för att tillmötesgå det portugisiska rådsordförandeskapet .
Likaså lägger ni vikt vid direktivet om ramvillkor för vattenförsörjningen .
Också gällande detta vill jag be er att helt enkelt godkänna ändringsförslagen som parlamentet skall anta i Bryssel i februari - då lär vi få en bred enighet .
En sak till : Ni har sagt att ni vill koppla samman miljöpolitiken med den fysiska planeringen .
På den punkten kan jag ge er mitt fulla stöd .
Ni har möjlighet att på regeringskonferensen se till att det nya fördraget innehåller en europeisk kompetens för den fysiska planeringen .
Därmed skulle ni med ens ha vunnit över oss på er sida ; men att ni verkligen genomför det tvivlar jag starkt på .
Jag kommer dock att ge er mitt stöd för det .
Som avslutning en sak till : jag ber er att i samband med områdena miljöpolitik och integration i andra politikområden tänka på att det kommer att finnas en skyldighet att göra detta , liksom att dokumentera det .
Var vänlig och meddela era kolleger i medlemsländerna det och se till att den befintliga lagstiftningen verkställs ; när det gäller miljölagstiftningen är så inte alltid fallet .
Om ni gör det så har ni kanske inte utlovat lika mycket som vissa andra , men i stället utfört ett ordentligt arbete - och därmed önskar jag er lycka till .
Herr talman , herr rådsordförande !
Från det rika kölrummet på skeppet med de femton roddarna , det portugisiska ordförandeskapets fantastiska fynd av den europeiska symbolen , låt mig inrikta mig på Europas digitala utmaning .
Den digitala revolutionen är enligt min mening först och främst en revolution i systemet och kulturen när det gäller distribution av varor och tjänster .
Detta innebär att vi måste ta ställning till tre konkreta frågor som finns med i programmet .
För det första tvingar den oss att på nytt reflektera över jämvikten mellan den offentliga och den privata lagstiftningen , jämvikten mellan lag och det som vi skulle kunna kalla soft law .
Anledningen är att - som någon sade vid Madridkonferensen - att ett år motsvarar två månader och fyra år , som är en skälig tid för handläggandet av ett normalt direktiv , motsvaras i det här fallet av 24 år .
En alltför lång tid .
För det andra måste vi väcka förtroende hos konsumenterna och de små och medelstora företagen samt skapa ett klimat och en kultur av kontrollerad risk , även om det kan verka motsägelsefullt .
För konsumenternas räkning måste vi sätta igång kommissionens utmärkta initiativ om en utomrättslig lösning av konflikter , som en följd av Tammerfors , men konsumenterna måste också betraktas som vuxna .
För de små och medelstora företagen måste vi förstärka den dialog som inletts med företag och konsumenter inom ramen för den inre marknaden .
Men även mera konkreta frågor , som till exempel att inta en fast ståndpunkt i enlighet med den affärsmässiga kulturen när det gäller artikel 15 i de nya Bryssel- och Luganokonventionerna , annars kan hela projektet om E-Europa gå i stöpet .
Avslutningsvis , och här sluter jag upp bakom Cox , så har vi utmaningen i den transatlantiska dialogen .
Inget är uträttat så länge som vi inte minskar avståndet mellan oss och Förenta staterna , dock i samordning med dem .
I den här frågan tror jag att vi behöver god samordning , ett bra samarbete och givetvis mycket uppmuntran .
" Skeppet seglar " - var de portugisiska styrmännens uppfattning på medeltiden .
Våra styrmän under de här sex månaderna är duktiga , det är jag övertygad om . )
Herr talman , ärade kollegor !
Jag har två för mig grundläggande frågor när det gäller det portugisiska ordförandeskapets ambitiösa halvårsprogram : det ekonomiska samarbetet med medelhavsländerna samt de främjande- och sysselsättningsbevarande åtgärderna .
Herr talman , parlamentet antog i november en resolution där man inom ramen för associeringsavtalet tog det alltmer intima samarbetet mellan Marocko och Europeiska unionen i försvar .
Det vore oförståeligt om samarbetet när det gäller fiske nu skulle vara mindre .
Fiskerisektorn , ärade kollegor , är en mycket skör sektor .
Katastrofen med Erika visade detta klart och tydligt .
Portugals sjöfartstraditioner och de utmärkta förbindelser man har med Marocko borde användas , herr talman , för att gjuta mera blod i de för närvarande stillastående förhandlingarna om det nya fiskeavtalet .
Fiskerisektorn är koncentrerad till Europas minst gynnade områden och där är man i stort behov av den .
Vi behöver en ekonomisk , social och territoriell framstegsvänlig politik så att behållningen av den nuvarande ekonomiska blomstringen inte går till den mer framgångsrika industriella sektorn .
Jag uppmanar det portugisiska ordförandeskapet att visa beslutsamhet och mod inför den här utmaningen .
Herr talman , herr rådsordförande , herr kommissionär !
Jag tänkte ta upp två saker .
Den ena gäller en sammankoppling av transportpolitik och regeringskonferensen .
Det har av många kollegor redan framförts att vi inte vill ha en regeringskonferens som enbart behandlar leftovers från Amsterdam , utan att vi i viss men inte överdriven mån vill se en omfattande diskussion av nya befogenheter vilka behövs för att bibehålla Europeiska gemenskapens funktionsduglighet .
Ni i det portugisiska rådsordförandeskapet kan här göra något av avgörande betydelse för den europeiska transportpolitiken och för säkerheten och miljön i Europa .
Ni kan genomföra det parlamentet fattade beslut om i november : upprättandet av ett enhetligt europeiskt kontrollsystem för flygsäkerheten är en central fråga som måste behandlas i Europeiska unionen , vilket kan ske genom att denna punkt sätts upp på regeringskonferensens dagordning .
Men vi vill förvisso inte centralisera allt .
De operativa befogenheterna bör stanna kvar hos medlemsländerna eller hos privata organisationer .
Men styrfunktionen måste få en enhetlig europeisk reglering .
Den nuvarande splittringen i luftfarten leder nämligen till dröjsmål , förseningar och risker för passagerarna samt till en mycket stor och onödig belastning på miljön .
Ett europeiskt mervärde torde i första hand stå att finna i ett enhetligt system för flygsäkerheten i Europa .
På marken finns den inre marknaden , men uppe i luften råder splittring .
Det kan inte fungera bra .
Vi i Europaparlamentet står därför fast vid vår ståndpunkt och det är min förhoppning , herr rådsordförande , att ni stöder detta .
Det andra som ni kan göra för miljön , ekonomin och transporter är att snabbt formulera en gemensam ståndpunkt beträffande järnvägspaketet .
I december lyckades det finländska ordförandeskapet övervinna motståndet från den franska regeringen mot att öppna järnvägstrafiken .
Nu har jag åter känslan av att det är en tidsfråga .
Här har ni i det portugisiska ordförandeskapet en stor chans om ni bara kan formulera den gemensamma ståndpunkten inom kort .
Vi väntar på er åtgärd .
Vi vill att godstransporterna läggs om från vägarna till järnvägarna .
Hjälp oss med det !
Herr talman , kolleger !
Jag skall ta upp en fråga som ligger det portugisiska ordförandeskapet nära hjärtat , nämligen Angola , ett land där ett inbördeskrig har pågått i tjugofem år och som i dag är världens största humanitära katastrof .
Vi vet vilka som ligger bakom att Lusaka-avtalet inte har kunnat genomföras - det är i första hand UNITA .
Därför har världen också infört sanktioner mot UNITA .
Det finns också risker för en regional spridning av denna konflikt genom att regeringstrupper har gått in i grannstater och att UNITA har förenat sig med väpnade grupper i andra länder .
Humanitärt , som sagt , är detta världens största humanitära katastrof med två miljoner internflyktingar och ett ohyggligt lidande på båda sidor .
Vi vill därför att Portugal , inte minst dess regering , med sin demokratiska , antikolonialistiska tradition också uttrycker för parlamentet vilka åtgärder man avser att vidta för att på detta sätt göra något som kan bidra till en lösning .
Det är endast en politisk lösning som kan ge fred och försoning i Angola .
Herr talman , herr kommissionär !
Ni skall veta , herr rådsordförande , att er vilja att föra en dialog med Europaparlamentet sågs med blida ögon här , vilket inte är överraskande om vi tänker på den portugisiska regeringens långa erfarenhet av dialog .
Vi iakttar ordförandeskapets mål - vilka vi erkänner är ambitiösa - och ser olika prioriteringar , många som innehåller dialog och många frågor som skall inledas eller fortskrida .
Det oroar oss att vi ser färre frågor som kommer att avslutas och mål som skall uppnås , men vi hoppas innerligt att ordförandeskapet blir ett gott ordförandeskap , för hela Europa , för Europas medborgare och för portugiserna .
För Europa , som vi hoppas kunna hjälpa med uppbyggnad och förstärkning , och i vilket alla känner sig representerade och identifierade , ett Europa som inte bara är för några få eller där de stora kväver de små .
För detta Europa är det också än en gång nödvändigt , vid en tidpunkt då man överväger fördragsändringar , att ett ordförandeskap som utövas av ett litet land inte därför behöver vara sämre eller mindre effektivt än det som utövas av de stora länderna .
För de europeiska medborgarna som vill ha ett Europa som engagerar sig i deras problem och inte bara i sina bankkonton eller sina produkter , som vill ha ett Europa som bryr sig om säkerheten , kampen mot droger och brottslighet , kontrollen av den illegala invandringen och antagandet av åtgärder för ett område med frihet , säkerhet och rättvisa .
Jag är säker på att ministern håller med mig i mitt positiva omdöme av den stora kompetens och kvalitet som den portugisiske kommissionären , António Vitorino , besitter och jag hoppas att rådet , i de områden han har fått hand om , kan ta konkreta steg enligt den scoreboard som beslutades i Tammerfors .
Och för portugiserna , som minns det goda ordförandeskapet för rådet när Portugal utövade det första gången för exakt åtta år sedan , och vi hoppas att den socialistiska regeringen kan leva upp till det prestigefyllda och effektiva arvet .
Herr talman , kära kolleger och herr rådsordförande !
Ni , herr rådsordförande , försöker skapa en mer positiv attityd till Europaparlamentet .
Ni accepterar de europeiska medborgarnas röst som en del i det europeiska beslutsfattandet , vilket vi uppskattar .
Vi hoppas och räknar med att denna positiva attityd håller genom hela sexmånadersperioden .
På rättsområdet är det nödvändigt med europeiska åtgärder .
Ni lyfter fram frågan om brottsoffer .
Det är en fråga som symboliserar medborgarnas rättssituation ur väldigt många dimensioner .
Det handlar om att inte längre diskriminera de medborgare som nyttjar sin fria rörlighet .
Jag har länge kämpat just för att förstärka brottsofferskyddet .
Om staterna inte är beredda att värna individerna och mildra våldets konsekvenser , så kan vi aldrig skapa den säkerhet som alla talar så vackert om .
Utan fördragsfästa , individuella medborgerliga rättigheter och tillräckliga resurser för polis och rättsväsende får vi inte den frihet och trygghet som medborgarna i Europa förväntar sig .
Ni kan driva på processen genom att öppet använda resultattavlan och visa att vi behöver framsteg .
Tidsgränser för åtgärderna skulle kunna öka takten .
Ni måste genomföra nödvändiga prioriteringar i ert ambitiösa program .
Då skulle jag vilja framhålla brottsoffer , scoreboard och organiserad brottslighet .
Jag hoppas att ni vill bekräfta att det är dessa frågor och medborgarrättigheterna som står allra överst på er prioriteringslista .
Därmed vill jag önska lycka till och stor framgång .
Det är glädjande att kunna konstatera att Afrika hör till det portugisiska ordförandeskapets prioriteter .
Europa har här verkligen ett stort historiskt ansvar och det skulle vara mycket oansvarigt att överlåta den svarta kontinenten till amerikanerna .
Jag hoppas att det euro-afrikanska toppmötet blir av och att unionen äntligen lyckas anta en gemensam ståndpunkt med avseende på konflikten i Centralafrika .
Det är logiskt att Portugals uppmärksamhet främst riktas mot Angola .
Jag vill ändå göra några randanmärkningar angående utlåtandet om kriget i Angola där rebellrörelsen UNITA utpekas som huvudskyldig .
Det är mycket riktigt så att Savimbi sköt sönder det första fredsavtalet när han förlorade valet 1992 .
Det är också lika riktigt att UNITA har använt avväpningsperioden till att beväpna sig igen och att de i det pågående kriget gjort sig skyldiga till grova kränkningar av de mänskliga rättigheterna .
Det måste vi fortsätta att fördöma .
Det gör dock inte att ledarna i Angola går fria .
Det var ju regeringen som i slutet av 1998 förklarade totalt krig mot rebellerna och som inte heller sparade civilbefolkningen i det kriget .
Det står också lika klart att även regeringen har beväpnat sig rejält under den här fredsperioden .
Människorättsorganisationer som Human Rights Watch och Global Witness anklagar regeringen för korruption i stor skala , för att använda miljarder oljedollar till militära inköp , bland annat från Portugal , och för förtryck mot oppositionen och mot pressen .
Afrikas näst största oljeproducerande land har en av de sämsta socialekonomiska indikatorerna i världen med undernärda barn och koleraepidemier ända in i huvudstadens centrum .
Europa måste fortsätta yrka för en dialog utan att gå in i en militär logik .
Portugal kan i det avseendet spela en viktig roll .
Inte genom att inta en ensidig hållning men genom att påpeka för båda parter det ansvar de har .
På det sättet kan det äntligen skina litet ljus i den mörka angolanska tunneln .
Herr talman , bästa företrädare för rådet !
För det första vill jag instämma i min kollega Coelhos ståndpunkt att ett litet land på ett märkbart sätt verkligen kan föra unionen framåt under sitt ordförandeskap .
Detta bevisade vi under det finländska ordförandeskapet , och jag är säker på att även Portugal kommer att lyckas med detta arbete .
Den kanske största utmaningen som Finland lämnade över till Portugal är slutförandet av det så kallade skattepaketet i samband med uppförandekoden för beskattning .
När Portugal för första gången redan före årsskiftet efter toppmötet i Helsingfors informerade de övriga medlemsstaterna om var man tänkte lägga tyngdpunkten under sitt ordförandeskap var jag synnerligen besviken på det sätt som man talade om skattepaketet , precis som om man redan hade avstått från försöken att uppnå en kompromisslösning .
Förra veckan uppträdde emellertid Ekofin-rådets nya ordförande Pina Moura på ett betydligt stramare sätt och återgav mig tron på att Portugal i likhet med det tidigare ordförandelandet Finland anser det viktigt att harmonisera beskattningen i medlemsstaterna på det sätt som föreslås i skattepaketet .
Det var också glädjande att höra att skattepaketet även i fortsättningen kommer att behandlas som en helhet .
Det är inte fråga om ett hopplöst fall .
Redan i resolutionen från toppmötet i Helsingfors kom medlemsstaterna överens om principen att alla unionsmedborgare skulle betala en lämplig skatt på alla inkomster från sina besparingar .
Denna lämpliga skatt kan förvisso utformas på många olika sätt .
Det är alltså viktigt att också rikta uppmärksamheten på olika typer av informationsskyldighet , detta för att säkerställa en rättvis och heltäckande beskattning .
Jag hoppas därför att rådet så snabbt som möjligt utser den skatteutredningsgrupp på hög nivå som var på tal redan i Helsingfors och fortsätter där man stannade i Helsingfors .
Utöver skattepaketet växer trycket på att åstadkomma ett enhetligt energiskattesystem som är neutralt i förhållande till det totala skattetrycket .
För egen del stöder jag varmt detta mål , om reformen bara genomförs utan att äventyra den europeiska industrins konkurrenskraft .
Den tredje utmaningen i fråga om beskattning är förknippad med mervärdesskatten .
Vårt mål är att övergå till ett slutgiltigt mervärdesskattesystem så snart detta är möjligt .
Jag hoppas att man håller även detta i minnet under den portugisiska perioden .
Herr talman !
Herr tjänstgörande rådordförande , ni har verkligen utarbetat ett ambitiöst verksamhetsprogram .
Vi i Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater gör oss stora förhoppningar om detta på det planerade toppmötet om sysselsättning .
De krav som den kristdemokratiske ministerpresidenten i Luxemburg Juncker formulerade inför sysselsättningsmötet 1997 omfattar också det planerade särskilda toppmötet i Lissabon .
Det får inte bara bli ett toppmöte på papperet , vilket varit fallet i otaliga icke bindande förklaringar på många toppmöten - Juncker pekade på det .
Däremot nådde regeringscheferna en konkret framgång med det så kallade Luxemburgförfarandet , dvs. en samordning genom sysselsättningspolitiska riktlinjer samt nationella handlingsplaner .
Sedan 1997 har dock de riktigt stora framgångarna låtit vänta på sig .
Det är framför allt när det gäller det praktiska genomförande av riktlinjerna som bristerna visar sig .
I det gemensamma sysselsättningsbetänkandet från 1999 räknas i detta sammanhang upp olika åtgärder som saknas i medlemsländerna ; det gäller reformen av skatte- och socialförsäkringssystemen , uppslutningen kring idén om livslångt lärande , brister i samband med främjandet av samarbetet mellan arbetsmarknadens parter med syftet att modernisera arbetsmarknadens struktur .
Sysselsättningspolitiken spelar sedan många år en viktig roll i parlamentet .
Men dessvärre har råd och regeringschefer knappt övertagit någonting av innehållet i våra förslag under 1999 heller , det gäller bland annat den så kallade europeiska sysselsättningspakten i Köln eller riktlinjerna 2000 .
Jag ber det portugisiska ordförandeskapet att göra vad det förutskickat i sitt PM för eftertanke : gör det bara ännu bättre och ta större hänsyn till vad vi säger !
En ny ekonomisk dynamik , konkurrens och flexibilitet måste bringas till överensstämmelse med de grundläggande behoven av social trygghet .
Den sociala marknadsekonomins framgångsrika princip är framtidsmodellen för Europa .
Ordförande Gama !
Vi uppskattade mycket det ni sade om parlamentets roll , om regeringskonferensen och om ledamotsstadgan , men vi måste också tala om utvidgningen av Europeiska unionen .
Utvidgningen österut är viktig , vi vill skapa ett politiskt Europa , men vi måste se till - och Portugal , precis som Italien är ett Medelhavsland - just när det gäller det stora Medelhavsområdet så att vi också skapar en välbehövlig Medelhavspolitik och balanserar utvecklingen österut mot en utveckling söderut .
När det gäller Europeiska rådet så tror jag att det är tre frågor som man måste diskutera .
Ni talade om sysselsättningen och för oss är detta utomordentligt viktigt , det är den allra viktigaste frågan .
Vi kämpar genom att hjälpa de små och medelstora företagen , få fart på turismen genom utvecklingspolitik och genom att kraftigt sänka skattetrycket .
Något annat som ligger oss varmt om hjärtat - det underströk ni själv - är frågan om rättssystemet .
Politiken när det gäller rättssystemet i Europa är mycket viktig .
Här förekommer alltför utdragna processer , felaktiga processer - och Italien har tyvärr ett negativt rekord i det avseendet - och även i flera av Europas länder ett politiserat rättssystem där vissa domare använder sin makt , inte för att utöva sina ämbeten , utan för att bedriva politik och ofta för att komma åt oppositionen och olika minoriteter .
Jag vill avslutningsvis peka på en tredje fråga efter sysselsättningen och rättsväsendet : narkotikaproblemet .
Detta är en viktig social fråga som vi känner särskilt starkt för , eftersom den berör miljontals ungdomar .
Kampen mot narkotikan borde vara en av det portugisiska ordförandeskapets , Europeiska kommissionens och detta parlaments viktigaste uppgifter .
Kampen måste föras mot de gamla , men även och framför allt mot de nya drogerna , utan att man faller för frestelsen att liberalisera drogerna , utan att man faller för frestelsen att legalisera och godkänna ett terapeutiskt bruk av ämnen som heroin , något som detta parlament redan har tillbakavisat .
Miljontals ungdomar följer oss uppmärksamt : de följer vad som sker i EU och av EU förväntar de sig ett svar .
Herr talman !
Jag skulle vilja göra tre kommentarer .
Den första gäller Sydosteuropa och Medelhavet .
Alla känner till att det är en orolig region , och den som trodde att problemen skulle kunna lösas under det portugisiska ordförandeskapets sex månader skulle vara naiv .
Jag uppmanar emellertid ordförandeskapet och kommissionen att göra allt vad som står i deras makt för att göra det möjligt för organisationen för Balkans återuppbyggnad , som har sitt säte i Thessaloniki , att på bästa möjliga sätt att uppfylla sitt uppdrag .
Jag skulle också önska , å ena sidan , att Turkiet inser att statusen som kandidatland medför skyldigheter att rätta sig efter gemenskapens regelverk och , å andra sidan , att ordförandeskapet och kommissionen påminner landet om dessa skyldigheter .
Min andra kommentar gäller regeringskonferensen .
Det skulle vara rätt att införliva stadgan om de mänskliga rättigheterna i det nya , reviderade fördragets text , för det är något som i mycket hög grad intresserar Europas medborgare .
Dessutom bör dagordningen utvidgas .
Det bör finnas en rättslig grund för en gemensam försvars- och utrikespolitik .
Särskilt vill jag påminna om en sak som parlamentet också har givit sitt stöd åt i betänkandet av Dimitrakopoulos-Leinen , det vill säga att det bör avsättas nya medel till viktiga och framträdande frågor , som till exempel turism och kultur .
Den tredje kommentaren gör jag i egenskap av ordförande i utskottet för regionalpolitik , transport och turism .
Ert program , herr rådsordförande , har rätt inriktning , men vi skulle förvänta oss att ni var mer optimistiska .
Jag skulle särskilt vilja understryka att det för oss är nödvändigt att frågan om åtgärdspaketet för avregleringen av järnvägarna avslutas under det portugisiska ordförandeskapet och att man arbetar för en lösning på problemet med förseningarna i luftfartssystemet .
Vi bör alltså övergå från dagens mellanstatliga system , Eurocontrol , till ett enhetligt system , där kommissionen bör ha initiativet , så att vi kan få ett slut på de hela tiden allt värre problemen för passagerarna som flyger över Europa .
Herr talman , herr rådsordförande , herr Costa , herr kommissionär !
Det är tydligt att det portugisiska ordförandeskapet har en mycket tung ansvarsbörda under de kommande sex månaderna .
Jag vill lyckönska ordförandeskapet när det gäller genomförandet av denna ansvarsbörda .
Prioriteringarna i sammanhanget riktas naturligtvis mot utvidgningen av Europeiska unionen - en utvidgning som i omfattning och karaktär skiljer sig från alla tidigare utvidgningar .
Vi vet också att EU : s utrikespolitik sträcker sig in i Östeuropa och att handlingsplanen för den gemensamma strategin i Ukraina redan gett resultat sedan toppmötet i Helsingfors , i och med tillkännagivandet om att dödsstraffet avskaffats .
I den inledande meningen i sitt tal till oss i förmiddags berörde utrikesminister Gama folkopinionens betydelse och hur viktigt det är att lugna medborgarna i Europeiska unionen .
Jag har bara en fråga som rådsordföranden kanske kan ta upp i sitt svar .
Kan han försäkra oss att hans oro rörande folkopinionen omfattar folkopinionen i ansökarländerna i Central- och Östeuropa ?
Han kanske inte anser att detta är en lämplig tidpunkt för att informera om vilka initiativ han har i åtanke för att se till att inte bara tempot i förhandlingarna upprätthålls , utan också att stöd till ansökarländerna säkerställs .
Jag skulle uppskatta ett lugnande svar från hans sida .
Herr talman !
Jag vill understryka ett par punkter som enligt min åsikt tas upp på ett mycket positivt sett i det portugisiska ordförandeskapets program .
Det gäller nödvändigheten att förena unionens utvidgning med institutionella reformer som kan garantera EU : s politiska roll , i enlighet med vad parlamentet har begärt av regeringskonferensen .
Europa har nu till sitt förfogande en inre marknad och en gemensam valuta .
Men trots detta är det nu dags att med större kraft ta itu med arbetslösheten och att åter börja driva frågan om en harmonisering av skattepolitiken och den sociala politiken , grundläggande faktorer i den sociala sammanhållningen .
Vi måste förstärka vår konkurrenskraft i en allt mer globaliserad ekonomi som har att möta utmaningen från informationsrevolutionen .
Här behövs en ny strategi för forskning , förnyelse och utbildning , frågor som det dokument som godkändes i går av kommissionen kommer att starta en viktig debatt om .
Utvidgningen av unionen , som i första hand vänder sig österut , är en verklighet och ett framtidsperspektiv som berör samtliga europeiska länder .
Jag håller emellertid med det portugisiska ordförandeskapet om att denna prioritering inte får minska uppmärksamheten gentemot Medelhavet , för fred och utveckling i det området är något som direkt berör Europas framtid .
Herr talman , mina damer och herrar !
Denna debatt har varit av alldeles särskild nytta för ordförandeskapet och vi kommer att med största uppmärksamhet ta till oss och analysera de förslag och anmärkningar som har lämnats här .
Under detta ordförandeskap kommer vi att arbeta mycket tillsammans med Europaparlamentet , även med kommissionen , den höge representanten Javier Solana och Västeuropeiska unionen , för vilken vi också är ordförandeland , och vi hoppas att detta samarbete kommer att bli fruktbart i hela ordets bemärkelse .
Vi bär med oss uppfattningen härifrån att det portugisiska ordförandeskapets grundläggande inriktning har ett enhälligt stöd och att det har bekräftats av Europaparlamentet , detta är viktigt för oss eftersom det stimulerar oss att arbeta i större samstämmighet .
När det gäller frågan om sysselsättning och innovation ser det extra toppmötet i Lissabon i parlamentet en extremt uppmärksam kammare , intresserad och engagerad i att göra Europa , under det sekel vi nu inleder , på samma gång till ett område med social sammanhållning och det mest dynamiska ekonomiska området i världen , för att möta globaliseringen och för att kunna demokratisera informationstekniken , och skapa en kunskapsekonomi , fri från mönstren och kännetecknen i en ren produktionsekonomi .
Även att genomföra utvidgningen , detta historiska tecken för slutet på det kalla kriget och bygget av det återförenade Europa .
Angående Turkietfrågan så skall vi noggrant fördjupa den för att samtidigt verka genom gemenskapens regelverk , screening , tillämpningen av Köpenhamnskriterierna och det strategiska målet att göra Turkiet till ett land med inriktning på att stadigt närma sig Europa .
Jag vet att detta parlament hyser vissa tvivel om detta .
Men jag skulle också vilja lugna er genom att säga att en annan politik skulle vara ännu värre för Europa , det skulle vara mycket negativt och få allvarliga konsekvenser för det vi vill med unionen , såväl internt som på ett internationellt plan .
Beträffande regeringskonferensen tycker jag att det har gått bra att få till en förtroendefull enighet mellan ordförandeskapet och parlamentet när det gäller behovet att integrera det senare på ett mer substantiellt , verkligt och kontinuerligt sätt i förhandlingsprocessen .
Och vi är öppna för detta .
I det brev jag skickade till parlamentets talman i början av det portugisiska ordförandeskapet gjorde jag till och med klart att vi , i egenskap av ordförandeskap , stod till förfogande för att delta i möten med ert utskott för konstitutionella frågor , och även i kammaren , om Europaparlamentets kammare en dag mer djupgående vill diskutera de ämnen som kommer att tas upp på regeringskonferensen .
Denna kommer att respektera maktdelningen , varje organs ansvarsområde , men jag tror att den kommer att stimulera den europeiska debatten om den institutionella reformen .
Det finns ingenting som hindrar oss från att agera på detta sätt .
Vi har för övrigt inte någon låst syn i förhållande till Helsingforsdagordningen .
Detta gör det möjligt , enligt de termer som formulerats , att införa vissa nya punkter .
Jag har själv diskuterat denna punkt med mina kolleger , i den rundresa jag gjorde till de europeiska huvudstäderna .
Statssekreteraren för Europafrågor kommer också att göra det nu .
Jag skrev till mina europeiska kolleger , till utrikesministrarna , i början av januari , för att be dem nämna de punkter de respektive regeringarna såg som möjliga att lägga till dagordningen för leftovers , så att vi mycket tidigt under ordförandeskapet och regeringskonferensen , skulle kunna få en tydlig bild av detta problem som vi också skulle kunna dela med Europaparlamentet .
Jag skrev även till kollegerna i ansökarländerna , både till dem i första och i andra utvidgningsomgången - vilka vi för övrigt hoppas skall kunna bli en enda linje - , för att be även dem att uttrycka sin åsikt om regeringskonferensen , för det värsta som kan inträffa när det gäller utvidgningen av Europa är att den institutionella reformen i Central- och Östeuropa skulle uppfattas som en slags förebyggande åtgärd mot dem som skall ansluta sig .
Det skulle skapa en relation full av misstroende .
De åtgärder som konferensen måste vidta är åtgärder för att få Europa att fungera bättre , det handlar inte om åtgärder för att förhindra anslutningsländerna att en dag kunna göra sin röst hörd inom det europeiska beslutssystemet .
Därför är det viktigt att de redan nu deltar och att vi lyssnar på deras åsikter .
Därför kan vi tycka att det inte är orealistiskt , som en av ledamöterna sade , att vi nu , under Europeiska rådet i Lissabon , försöker få en tydligare bild , om vi är överens om vilket spektrum vi kommer att ha , av regeringskonferensens dagordning .
När det gäller den gemensamma säkerhets- och försvarspolitiken handlar det om en dimension som saknas för att kunna hävda Europa på ett utrikesplan .
Europeiska unionens utrikespolitik kommer inte att vara någonting så länge den inte innehåller denna komponent .
Vi kommer under detta halvår att ta avgörande steg för att denna skall kunna skapas , vi kommer att genomföra den första övning där Nato överför kapacitet till Västeuropeiska unionen och denna kommer att verka under Europeiska unionens politiska riktlinjer .
Men var lugna , kolleger och ledamöter från medlemsstater som är medlemmar i Atlantpakten : denna övning kommer att genomföras inte för att minska utan för att öka den europeiska säkerheten .
Detta innebär hela tiden en mycket uppmärksam och mycket omdömesgill relation till dem bland oss som inte är med i Atlantpakten , men som kan få tillgång till alla dessa system om de önskar .
Och om de vill detta , kommer de att medverka på jämlik grund med övriga partner .
Angående några punkter i utrikespolitiken som ledamöterna tog upp , när det gäller toppmötet Europeiska unionen / Afrika : vi har inte med detta som ett uttryckligt mål för det portugisiska ordförandeskapet , när vi tog emot ordförandeskapet ansåg vi att detta mål inte var tillräckligt klart och vi ville inte göra européerna besvikna genom att införa en ram som vi inte hade några garantier för .
Vår arbetsordning är följande : vi fortsätter att arbeta för att när som helst kunna återuppta denna idé , om det är möjligt att göra det i tid och under logistiska villkor för att kunna genomföras .
I annat fall kommer vi att fortsätta att fördjupa dess behandling tillsammans med våra afrikanska partner , och vi kommer att skapa en grund för att detta skall kunna tas upp och genomföras i framtiden .
Problemet med vapenembargot mot Indonesien : i september , under det mest dramatiska ögonblicket i Östtimors drama , beslutade Europeiska unionen att för en begränsad period , vilken upphör nu i januari , införa ett vapenembargo mot Indonesien .
Den lösningen innehöll ingen mekanism för en automatisk förlängning och möjligheten att uppnå enhällighet i rådet var att nu inte lägga fram något nytt vapenembargo mot Indonesien , utan att med all tydlighet understryka att Europeiska unionens medlemsstater i denna mening är underställda en sträng uppförandekod som innebär mycket stränga regler för slutdestinationen av vapnen och för dess användning .
Vårt enhälliga beslut var mycket tydligt när vi betonade att denna fråga fortsättningsvis kommer att vara föremål för granskning och att embargot är en mekanism som Europeiska unionen när som helst kan ta till , så som den har gjort , för att ingripa och använda sig av i dramatiska situationer för att lösa dessa och hejda dem .
När det gäller Angola handlar det om ett land med oerhörda resurser och med en sällsynt egenskap i Afrika , att inte bestå av en omåttligt stor befolkning , varken i förhållande till landets storlek eller till sina resurser .
Angola har dragits med en konflikt , en osäker situation , och lider också av stor livsmedelsbrist och stora humanitära problem .
Lusakaavtalen har inte uppfyllts av en av parterna .
En av de viktigaste frågorna i den angolanska processen har varit att en av parterna har vägrat avmilitarisera sig för att övergå till att bli ett civilt parti som kan ingå i ett normalt institutionellt system .
Det är viktigt att detta sker och därför är Europeiska unionens beslut inriktat på att stimulera alla de som i ett av områdena , UNITA : s , vill och är beredda att verka på politisk väg och inte genom vapen .
Men det finns också behov som alla erkänner .
Jag var i Angola för omkring fyra dagar sedan och jag talade inte enbart med presidenten och regeringsmedlemmarna , utan också med ledamöter från alla parlamentariska riktningar , även de ledamöter som vi kan räkna till UNITA : s olika tendenser , och jag kunde dra slutsatsen att ett stort antal anser att en förbättring av det angolanska systemet är nödvändig .
Några av dessa förbättringar håller på att inledas och det är nödvändigt att stimulera deras förverkligande : en förbättring av det finansiella systemet , en förbättring av landets nationalräkenskaper , av insynen i dem och deras bestämmelser .
I detta syfte kommer säkert inledningen av förhandlingarna med Internationella valutafonden och ett eventuellt undertecknande av en första överenskommelse , inom kort att skapa lämpliga förutsättningar för att inom ramen för Parisklubben kunna utforma en bilateral mekanism för att övervaka regleringen av Angolas skuld , vilket gör det möjligt för Europeiska unionen att lösgöra de medel som beslutades för flera år sedan , under rundabordskonferensen om Angola , men som än i dag hålls inne av de skäl vi känner till .
En förbättring av det institutionella systemet , med en konstitutionell revidering vars debatt naturligtvis inleds med antagandet av de pluralistiska värdena , rättsstaten och pressfriheten .
Jag vill här betona betydelsen av den debatt som kommer att äga rum i det angolanska parlamentet om journalisternas rättigheter och det grundläggande behovet av en oberoende press i ett modernt politiskt system .
Det är uppenbart att detta kommer att gagna en återvändo av Angola till det internationella systemet , en förbättring av FN : s eget system , vilket är extremt viktigt .
Jag vill därför framhäva det faktum att förhandlingarna mellan den angolanska regeringen och FN : s generalsekreterare har lett till ett öppnande av ett FN-kontor i Angola med övervakningsfunktioner och arbete med humanitär hjälp , vilket kommer att få stor betydelse för den angolanska befolkningen .
Det krävs således , samtidigt med den nödvändiga avmilitariseringen av ett politiskt parti , en institutionell förbättring , en förbättring av det finansiella systemet och av systemet för samordning med FN-organisationernas allmänna ram .
Europeiska unionens medverkan i denna process är givetvis av stor betydelse , dels för den omedelbara humanitära hjälpen , dels för utarbetandet av ett stödprogram till återuppbyggnad och återanpassning .
Herr talman , ärade ledamöter !
Det är omöjligt för mig , av tidsskäl och genom att en ny punkt om Mellanöstern tillkommit i er arbetsordning , att förlänga mitt anförande mer , men jag skulle vilja avsluta med att säga att det är mycket tillfredsställande för ordförandeskapet att här i debatten se hur vi kan uppnå en allmän samstämmighet om våra föreslagna grundtankar och även att det var möjligt - vilket jag också tycker att vi har uppnått - att definiera en arbetsmetod med Europaparlamentet som jag är säker på kommer att bidra till att berika rådet och Europaparlamentet inom den allmänna verksamhetsramen för våra institutioner .
( Ihållande applåder ) Tack så mycket , herr rådsordförande .
Jag förklarar debatten avslutad .
 
Fredsprocessen i Mellanöstern Nästa punkt på föredragningslistan är rådets och kommissionens uttalanden om fredsprocessen i Mellanöstern .
Herr talman , mina damer och herrar !
Jag skall mycket kortfattat säga att jag precis har kommit tillbaka , med höge representanten för den gemensamma utrikes- och säkerhetspolitiken , Javier Solana , med Europeiska unionens specielle sändebud , Miguel Moratinos och med representanten för en av kommissionärerna , från en resa till Mellanöstern , där vi för unionens räkning fick träffa de högst uppsatta personerna i Syrien , Israel , de palestinska områdena , Jordanien , Egypten och Libanon , och vi hade även ett möte med generalsekreteraren för Arabförbundet .
Fredsprocessen i Mellanöstern har en god inriktning , på ett allmänt plan , men den möter två omedelbara flaskhalsar : en är den israelisk-palestinska komponenten , som gäller vissa förseningar i tidsplaneringen och även det uppskjutna datumet för förhandlingsstarten av slutstadgan , den andra handlar om den syriska sidan , med förseningar på grund av Syriens vägran att tillfälligt fortsätta förhandlingarna i Washington .
Denna försening av den syriska frågan har stor betydelse , då den försvårar och villkorar inledningen av förhandlingarna om Libanon .
Europeiska unionen har genom åren bedrivit ett mycket konsekvent progressivt arbete genom det speciella sändebudet Miguel Moratinos , vars arbete jag vill betona , genom ett kontinuerligt arbete av kommissionen och nu av den höge representanten ; och detta besök kommer att få sin fortsättning då president Arafat , på måndag , besöker rådet ( allmänna frågor ) , efter sin resa till Washington , och liksom vi redan har träffat Israels utrikesminister Levy , planerar vi inom kort ett möte med Syriens utrikesminister inom ramen för de fortsatta förhandlingarna .
Vi kommer också att delta - ordförandeskapet , kommissionär Christopher Patten och den höge representanten - i det multilaterala mötet i Moskva den 1 februari , där vi kommer att lägga fram Europeiska unionens ståndpunkter .
Unionen har , utan att vara part i förhandlingarna , ständigt arbetat för att stödja och befästa fredsprocessen , med stark närvaro i den multilaterala processen och får i februari tillfälle att åter sätta i gång arbetet i arbetsgruppen om ekonomisk och regional utveckling som leds av unionen ; och vi har naturligtvis varit närvarande genom EU : s partnerskap med Medelhavsländerna i utarbetandet av en samling associeringsavtal med länderna i regionen , och ekonomiska biståndsprogram , och vi har även haft en närvaro genom Europeiska investeringsbanken .
Det finns ett medvetande i alla länder - detta kunde vi också konstatera under vår rundresa - , om att unionen , även om vi inte är part i förhandlingarna , men genom att vi är den viktigaste handelspartnern för praktiskt taget alla länder i området och den största givaren av offentligt stöd till de palestinska områdena , på medellång och lång sikt har en oumbärlig roll att spela i att etablera fred i Mellanöstern , och det finns redan nu lämpliga ramar som utvecklas för att ge verklig form åt detta samarbete , dels i flyktinghjälp , dels i utarbetandet av integrerade samarbetsprogram , främst för att lösa vattenproblemet , både för hela vattenhanteringen , och vad gäller specifika regionala utvecklingsprogram .
Det var också möjligt att se till att vår medverkan i denna process inte skedde i motsättning till USA , utan genom ett regelbundet meningsutbyte och vårt uppdrag , som slutade i går , ledde till slutsatsen att det behövs en förstärkning av unionens redan stora engagemang i hela Mellanösternfrågan .
Detta är ännu en punkt där det är absolut nödvändigt att ha ett ständigt samarbete mellan rådet och kommissionen , och även ett ständigt samarbete mellan dessa två organ och parlamentet .
( Applåder ) Tack så mycket , herr rådsordförande , för ert uttalande .
Vi avbryter debatten här för att inleda omröstningen .
 
OMRÖSTNING .
( NL ) Fru talman !
Jag ville bara göra mina tyska kolleger uppmärksamma på att det insmugit sig ett översättningsfel i en gammal version och jag vet inte om det har rättats till än .
Det gäller punkt 5 .
Där handlar det om budgetåret 1999 .
I den gamla tyska versionen står det 1997 .
Jag skulle också vilja klargöra , och jag har inte sett den senaste tyska versionen , att texten skall lyda på följande sätt : " förklarar att det inte kommer att vara berett att avsluta räkenskaperna för budgetåret 1999 om kommissionen inte åtgärdat de bokföringsfel som revisionsrätten påtalat " .
( Genom omröstning antog parlamentet i tur och ordning de två besluten och resolutionen . )
Betänkande ( A5-0001 / 2000 ) av van Hulten för budgetkontrollutskottet om åtgärder att vidta med anledning av den oberoende expertkommitténs andra rapport om reformering av kommissionen Beträffande punkt 48 Fru talman , jag har en begäran : i nästa punkt 48 handlar det om det känsliga ämnet kommissionärernas partitillhörighet .
På grund av att omröstningen om den första och andra delen kan missförstås eftersom det inte är fråga om någon första och andra del utan om en mellansats vi skall komma fram till , begär jag att ni läser upp mellansatsen så att samtliga kolleger vet vad de röstar om i dag .
Vi skall göra så här .
Beträffande ändringsförslag 27 Fru talman , ändringsförslag 27 är inte längre aktuellt då vi nådigt har fattat beslut om att vi faktiskt får bestämma våra egna regler , att vi bara tar råd från andra och att det inte är något annat organ som beslutar för oss .
De motsvarande orden har vi strukit och då har inskottet som skall läggas till med ändringsförslag 27 inte längre någon betydelse .
Det har bara en betydelse om ett annat organ beslutar om våra regler som det sedan kommer överens med oss om .
Men eftersom parlamentet har visat så pass ryggrad att det i vart fall gör anspråk på att bestämma över sina egna förfaranden så anser jag att ändringsförslaget inte längre gäller .
( Applåder ) Fru talman !
För tillfället kan jag inte hålla med föregående talare , eftersom detta har att göra med ledamotsstadgan .
Detta är skillnaden mellan parlamentet och rådet i detta fall .
Det är en helt annan fråga än den vi behandlade innan .
Vi står fast vid vårt ändringsförslag . .
( EN ) Fru talman !
Jag håller med Elles om att detta är en separat fråga , men jag håller också med Kuhne om att vi bör göra oss av med den .
Beträffande punkt 56 , ändringsförslag 6 .
( EN ) Fru talman !
Ändringsförslag 6 , i dess lydelse här , återspeglar inte på ett korrekt sätt den omröstning som hölls i budgetkontrollutskottet .
Jag har tagit upp saken med utskottets ordförande , som inte håller med om detta .
Men det är viktigt att framhålla här .
Låt mig förklara skillnaden .
Budgetkontrollutskottet röstade för den första delen av ändringsförslaget från utskottet för rättsliga frågor och den inre marknaden- eftersom det är vad detta är - och emot den andra delen .
Texten skall alltså lyda enligt följande : " ... anser att även om det totala löne- och förmånspaketet för tjänstemän måste vara attraktivt och konkurrenskraftigt när det gäller den övergripande nivån för ersättningar , behöver paketets struktur moderniseras . "
Utskottet föredrog den första delen , vilken är en språklig ändring , men var emot den andra delen , vilken är en innehållsmässig ändring .
Jag är rädd för att det är lite oklart för några av oss .
Alla har förstått er .
För min del låter jag det som står i texten gå till omröstning .
Fru talman !
Mellan den första och den sista versionen har Theatos betänkande om skydd för gemenskapens ekonomiska intressen genomgått en intressant utveckling .
Förslaget med en gemenskapsförordning om att inrätta en oberoende europeisk åklagare har fördömts , eftersom det uppenbarligen strider mot artikel 280 i fördraget , och har i stället omvandlats till en enkel uppmaning till den kommande regeringskonferensen .
Den har ersatts med förslaget om en förordning om att inrätta en ny ganska underlig enhet , en oberoende europeisk organisation som skulle kontrollera att de undersökningar som utförs av byrån för bedrägeribekämpning , OLAF , genomförs korrekt .
I detta andra förslag hittar jag på nytt mitt inlägg av den 25 oktober förra året , där jag liksom några andra parlamentsledamöter oroade mig över hur det interinstitutionella avtalet om OLAF : s undersökningar skulle tillämpas i Europaparlamentet .
Kanske man försöker att överväga vår kritik , även om det sker sent .
Tyvärr förefaller mig denna nya oberoende organisation som skulle kontrollera en oberoende byrå mycket underlig , och den besvarar fortfarande inte den grundläggande fråga jag ställde , nämligen vår kammares oberoende .
När det gäller den europeiska oberoende åklagaren är det ett förslag tvärtemot vår uppfattning om ett nationernas Europa , såsom jag förklarade i gårdagens debatt och i den debatt som ägde rum den 13 september förra året , om den andra rapporten från den oberoende expertkommittén .
En rad s.k. intellektuellt oberoende jurister fortsätter emellertid att lägga fram förslaget , men i verkligheten är de oftast betalda direkt eller indirekt av kommissionen , som enligt rapporten från den oberoende expertkommittén själv motarbetar kampen mot bedrägerier .
Vi finner det för övrigt otroligt att idén om en europeisk åklagare finns med i Theatos betänkande utan att man alls rådfrågat utskottet som ansvarar för att följa upp konstitutionella frågor , när en sådan innovation skulle ändra balansen mellan institutionerna på ett grundläggande sätt .
Men som vanligt när det gäller europeiska ärenden inleder man reformer utan att verkligen från början förklara hur omfattande effekterna blir .
Det ingår i den desinformation som gör att systemet fortsätter att fungera .
Fru talman !
Som företrädare för Pensionärspartiet röstade jag för förslaget att inrätta ett rättsligt skydd för unionens ekonomiska intressen .
Detta är och måste vara ett första steg mot skapandet av ett verkligt europeiskt rättsligt samarbetsområde när det gäller såväl civil- som straffrätt .
I annat fall hade jag inte röstat för förslaget , för det ligger inte i Europas intresse att inrätta ett rättsligt europeiskt organ enbart för att komma åt de egna bedrägliga anställda , de svarta får som det finns överallt .
Jag hoppas och yrkar på att medborgarna i hela Europa verkligen skall få en europeisk civilrätt och en europeisk straffrätt . .
( DA ) Vi har i dag röstat emot ett inrättande av ett europeiskt offentligt åklagarämbete av följande skäl : Vi stöder inte en gemensam europeisk straffrätt eller -myndighet .
Som utgångspunkt menar vi att man kan bekämpa kriminalitet lika effektivt med befintliga instrument , t.ex.
Europol och konventionerna om utlämning och inbördes rättshjälp .
I realiteten är det inte så stor skillnad mellan medlemsstaternas straffrätt att denna inte skulle kunna övervinnas med hjälp av de befintliga mellanstatliga instrumenten .
Vi kan emellertid fullständigt ansluta oss till kritiken av de 10 medlemsstater som ännu inte har ratificerat bedrägerikonventionen från 1995 .
Vi menar att det inte finns någon rättslig grund i fördraget för inrättande av ett europeiskt offentligt åklagarämbete .
Det finns inte stöd för att införa en myndighet som sysslar med frågor som berör medlemsstaternas straffrätt eller rättskipningsbestämmelser .
Ett alternativ till en europeisk offentlig åklagare skulle i stället kunna vara Eurojust , som föreslagits på toppmötet i Tammerfors .
En samordnande enhet bestående av nationella offentliga åklagare som skall stödja forskningen om brottsfrågor .
Vi välkomnar detta initiativ .
Det är precis ett sådant praktiskt samarbete det finns behov av .
Den europeiska offentliga åklagaren skulle först och främst bara kunna syssla med brott som begåtts av EU-anställda .
I realiteten finns det mer behov av en grundläggande reform av tjänsteföreskrifterna och de disciplinära förfarandena .
Det är bara de grövsta fallen som kommer att få straffrättsliga konsekvenser .
90 procent av fallen kommer att vara av disciplinär natur , som t.ex. försummelse eller inkompetens .
Det finns i stället behov av ordentliga interna kontrollförfaranden och en granskning av immuniteten för de anställda . .
( EN ) Låt mig säga när jag nu uttalar mig på den konservativa gruppens vägnar i Europaparlamentet , att vi betonar vårt engagemang när det gäller skyddet av Europeiska gemenskapernas ekonomiska intresse .
Vi skulle önska att konventionen och de två protokollen i detta sammanhang kunde undertecknas så snart som möjligt av alla medlemsstater .
Vi anser att det bör vara ett nära samarbete mellan medlemsstaterna för att se till att detta mål uppnås .
Men vi stöder inte idén om en enhetligt straffrättslig ram för att skydda EU : s ekonomiska intressen eller inrättandet av ett offentligt åklagarämbete på gemenskapsnivå .
Vi har därför i dag röstat emot Theatos betänkande .
Vi i frihetspartiet är ju sedan länge för effektiv kontroll och bedrägeribekämpning särskilt i samband med oegentligheter i EU : s budget .
Det är också grunden till vårt principiella gillande av Theatos betänkande .
Inte desto mindre är vi medvetna om framför allt den behörighetsrättsliga problematiken .
Mot bakgrund av detta uppmanas medlemsländerna att inom ramen för diskussionen om en reform av fördragen på nytt ta ställning till huruvida skapandet av egna EU-regler överhuvudtaget är meningsfullt och kommer att leda till målet .
Att det nuvarande rättsläget enligt vår uppfattning ej tolererar detta kan vi slå fast .
Den roll en " europeisk åklagare " - eller vad den än kallas - skulle få , skulle innebära allvarliga ingrepp i staternas suveränitet och kräver därför en grundlig diskussion .
Det förhållandet att bara ett fåtal medlemsländer har ratificerat avtalet om skydd för unionens finansiella intressen visar på nytt att möjligheterna för integrationen är begränsade .
Vi vill med bestämdhet understryka att en överföring av detta område till gemenskapen inte kommer i fråga och att en harmonisering av reglerna för brottsliga gärningar bör begränsas till de föreslagna områdena .
Skapandet av en enhetlig europeisk straffrätt motsvarar i vart fall inte våra föreställningar om i vilken riktning unionen bör utvecklas . .
( EN ) Detta betänkande handlar om skydd av Europeiska unionens ekonomiska intressen .
Det har visat sig att de metoder som för närvarande finns tillgängliga för att åtala personer som gjort sig skyldiga till bedrägeri i samband med EU-medel är olämpliga .
Det är t.ex. bara fem medlemsstater som ratificerat konventionen om skydd av Europeiska unionens ekonomiska intressen , trots att det passerat mer än fem år sedan de åtog sig att göra detta .
Den konservativa regeringen undertecknade inte konventionen , men labourregeringen följde nyligen Tysklands , Österrikes , Finlands och Sveriges exempel och undertecknade konventionen .
Under veckan när kommissionen sammanfattade sina reformförslag och betonade behovet av att förändra kulturen inom kommissionen , rekommenderade EPLP-gruppen genom sitt sätt att rösta , att tjänstemän som gjort sig skyldiga till överträdelser av gemenskapens bestämmelser skall åtalas .
Det nuvarande systemet för åtal mot tjänstemän som gjort sig skyldiga till överträdelser av gemenskapens bestämmelser fungerar inte , och detta är skälet till varför vi stöder uppfattningen om att ett offentligt åklagarämbete skall inrättas på gemenskapsnivå endast för personer som arbetar inom EU : s institutioner .
Vi har tydligt röstat emot alla förslag i sammanhanget som sträcker sig längre än så , och vi har kategoriskt röstat emot alla hänvisningar till Corpus Juris .
Genom vårt sätt att rösta har vi visat att EPLP-gruppen inte kan acceptera bedrägerier inom EU : s institutioner , och utmanar andra som har röstat emot detta betänkande att förklara hur de har tänkt sig att vinna kampen mot bedrägeri inom EU : s institutioner .
Betänkande ( A5-0004 / 2000 ) av van der Laan Fru talman !
I det betänkande som i dag lagts fram för oss föreslås att vi genom tillämpning av artikel 276 i fördraget skall bevilja kommissionen ansvarsfrihet för genomförande av Europeiska gemenskapernas allmänna budget för budgetåret 1997 .
De franska ledamöterna i Gruppen Unionen för nationernas Europa har vägrat att rösta för en sådan åtgärd .
Betänkandet om ansvarsfrihet för budgetåret 1997 ajournerades faktiskt av parlamentet redan den 4 maj förra året , eftersom det visade sig att Santers avgående kommission , som endast skulle sköta pågående ärenden , inte kunde göra åtaganden om reformer på sikt som föreföll nödvändiga , med tanke på den omfattande kritiken från revisionsrätten .
I dag har Prodis kommission åtagit sig detta och redan inlett flera reformer .
Men betyder det att vi skall bevilja ansvarsfrihet ?
Vi måste komma ihåg att revisionsrättens rapport om budgetåret 1997 var mycket sträng och man vägrade att bevilja någon revisionsförklaring om tillförlitligheten i de oegentliga transaktionerna enligt artikel 248 i fördraget .
Samtidigt som revisionsrätten nämnde att åtagandena föreföll riktiga lade den ändå till denna grundläggande precisering : " liksom tidigare år är inverkan av felaktigheterna i de oegentliga transaktionerna bland kommissionens betalningar av en sådan omfattning att revisionsrätten inte kan garantera att dessa transaktioner är lagliga och i sin ordning " .
Men om revisionsrätten inte vill avlämna sin revisionsförklaring om hela budgeten för år 1997 varför har då ledamöterna i Europaparlamentet beslutat att moraliskt godkänna den , genom att bevilja ansvarsfrihet ?
Naturligtvis invänder man att det inte handlar om samma kommission , men då svarar vi att genomförandet av budgeten för 1997 fortfarande är som det är .
Det har inte ändrats de senaste sex månaderna .
De oegentliga transaktionerna faller inte alla under kommissionens ansvar .
Medlemsstaterna har ofta också varit inblandade .
Fru talman !
För Pensionärspartiets räkning röstade jag för att kommissionen skulle beviljas ansvarsfrihet för budgetåret 1997 .
Men vad har pensionärer med ansvarsfriheten att göra ?
Jag minns att jag även har varit kamrer , och som sådan skulle det glädja mig om det kunde finnas så många euro som möjligt i de europeiska medborgarnas fickor .
Parlamentets kontroll när det gäller att bevilja ansvarsfrihet är med andra ord en viktig funktion och jag hoppas att såväl revisionsrätten som detta parlament skall få utökade befogenheter och framför allt att de skall få större möjligheter att utöva denna sin kontrollfunktion .
Jag skulle också önska att man var försiktig så att man inte spenderade tio euro för att de europeiska medborgarna skall få en .
Jag skulle dessutom önska att man garanterade en verksamhet som inte bara var formellt korrekt , utan som även var korrekt till sitt innehåll och i sin konkreta tillämpning .
Betänkande ( A5-0001 / 2000 ) av van Hulten Fru talman !
Van Hultens betänkande om reformerna avsedda att lösa kommissionens kris följer ganska troget den andra rapporten från den oberoende expertgruppen , som min grupp redan uttalade sig om den 13 september förra året .
Men de föreslagna reformerna sätts inte tillräckligt i sitt sammanhang , och det stora antalet förslag till punktförbättringar , ibland bra , ibland dåliga , kanske därför döljer de verkliga funktionsproblemen i de europeiska institutionerna .
Eftersom den första rapporten från den oberoende expertgruppen påvisade fall av individuella brister kunde man ha väntat sig att den andra analyserar korruption som förekommer permanent kring de europeiska institutionerna , såsom beskrevs i vissa dokument som cirkulerade i samband med att rapporten skrevs .
Men här finns inget av detta .
Det är naturligtvis bättre att föreslå framtidsreformer än att hela tiden gå tillbaka till det förgångna .
Men jag tror att dåtiden förbleknar och hindrar oss från att se omfattningen av de nödvändiga reformerna .
Dessa reformer är naturligtvis många , men vad det framför allt handlar om är frågan om kommissionens oberoende som förhindrar att man blir medveten om att den bara skall vara en enkel gemensam enhet för staterna , och som hindrar medlemsstaterna från att utöva en verklig kontroll över den .
Vi måste därför bekämpa allt som bidrar till att göra kommissionen till ett ogenomträngligt fort och bl.a. på nytt ge rådet en verklig politisk kontroll över kommissionen , stärka samarbetet i båda riktningarna mellan revisionsrätten och motsvarande nationella myndigheter för att förbättra kontrollerna både i staterna och i Bryssel , avskaffa de närmast diplomatiska privilegier som kommissionen åtnjuter och som motarbetar undersökningarna och öppna den europeiska offentliga funktionen mycket mer för nationella specialister på tillfälligt uppdrag .
Slutligen bör vi , såsom föreslagits av utskottet för sysselsättning och sociala frågor , i ett yttrande som inte resulterade i någon åtgärd , på nytt fullständigt se över möjligheten att finansiera intressegrupper , utan tillstånd i förväg , ur del A i budgeten , en möjlighet som i dag öppnar dörren för att dela ut anslag utan rättslig grund och gynnar klientilismen kring kommissionen .
Fru talman !
Som företrädare för Pensionärspartiet röstade jag för betänkandet om att reformera kommissionen .
I inledningen sägs det att vi röstar om denna förordning för att det är viktigt att återupprätta de europeiska medborgarnas förtroende för den europeiska integrationsprocessen .
Det är med andra ord rätt att det inte får förekomma bedrägerier och att det finns ett reglemente för kommissionen som skyddar oss mot risken att åter hamna i dessa situationer som , vilket jag redan påpekat , skulle kunna utgöra det enda svarta fåret .
Berthu , som talade före mig , har rätt : det som är viktigt är innehåller i det man gör .
Medborgarnas , och även de europeiska pensionärernas , förtroende uppnår man inte med hjälp av hundratusen förordningar och kommatecken utan framför allt med konkreta och kraftfulla handlingar från kommissionens sida , genom en minskning av antalet anställda i parlamentet , kommissionen och rådet . .
( DA ) Vi har i dag röstat för van Hulten-betänkandet , eftersom det innehåller många bra rekommendationer till reformering av kommissionen .
Vi vill särskilt lyfta fram en genomgripande reformering av personalpolitiken och en effektivisering och decentralisering av finanskontrollen .
Det finns emellertid enskilda punkter där vi har valt att rösta emot de framlagda förslagen .
Vi har röstat emot ett inrättande av en europeisk offentlig åklagare .
Vi menar att ett utvidgat mellanstatligt samarbete om forskning i brottmål , som föreslagits på toppmötet i Tammerfors , är en bättre idé .
Det finns dessutom snarare behov av en reformering av tjänsteföreskrifterna , eftersom bara ett fåtal fall får straffrättsliga konsekvenser .
Vi har röstat emot ett fullständigt avskaffande av förhandskontrollen .
Man skall behålla en viss förhandskontroll .
Det räcker inte med att bara ha en stickprovskontroll när pengarna betalats ut .
Man skall istället reformera och decentralisera kontrollen .
Vi har röstat emot en begränsning av parlamentets tillgång till information .
Parlamentet bör ha rätt till allt det material som kommissionen lämnade ut till den oberoende expertkommittén .
Vi har också röstat emot inrättandet av flera s.k. expertkommittéer .
Det bör vara de behöriga utskotten i parlamentet som genomför undersökningar och lägger fram förslag till reformer .
Faran med expertkommittéer är att man kan undergräva parlamentets roll som folkvald institution . .
( EN ) Herr talman !
Jag stöder helhjärtat min labourkollega Neil Kinnocks fina initiativ när det gäller att städa upp i den röra som Europeiska kommissionen lämnade efter sig .
På samma sätt som kommissionen inte kunde fungera med hjälp av teknik från 1950-talet , kan den inte heller fortsätta att fungera med en ledningskultur som praktiserades på 1950-talet .
Det finns ett desperat behov av en övergripande reformering av dess kontrollsystem för ledning och ekonomi .
Målet måste vara att skapa en effektiv , ansvarig och öppen kommission som medborgarna i Europeiska unionen återigen kan känna förtroende för .
Kommissionär Kinnock har fått en flygande start .
När det gäller att sortera bort obstinata , ålderdomliga organisationer som fastnat i sina dogmer , kan ingen jämföra sig med honom .
Hans förslag till en uppförandekod för alla tjänstemän inom kommissionen , avlägsnandet av nationell öronmärkning för höga tjänster och moderniseringen av förbindelserna med industrin är djärva , omstörtande och ett gott exempel på gammalt fint brittiskt sunt förnuft .
Det är faktiskt så att han tillför ett distinkt brittiskt drag av friska tag , effektivitet och ansvarighet till organisationen .
Det var naturligtvis Europaparlamentet och , framför allt , den socialdemokratiska gruppen under ledning av min f.d. kollega Pauline Green som tvingade kommissionen att öppna sig och erkänna att den behövde förändra sitt beteende .
Men vi kan inte slappna av riktigt ännu .
Kommissionär Kinnock har mött och kommer att fortsätta möta ett avsevärt motstånd mot reformerna .
Samtidigt som alla offentligt hävdar att de stöder en övergripande reform , finns det vissa eurokrater som egentligen gör vad som helst för att skydda sina hävdvunna intressen .
Inte heller de EU-fientliga från torypartiet kommer att missa några tillfällen då de kan vinna politiska poäng , inte ens på bekostnad av de mycket behövliga reformerna .
Brittiska ledamöter från den socialdemokratiska gruppen vid Europaparlamentet kommer emellertid även i fortsättningen att ge kommissionär Kinnock och hans reformprogram sitt fulla stöd .
Reformeringen får inte tappa fart p.g.a. själviska dagordningar som ställs upp av ett fåtal eurokrater och euroskeptiker . .
( EN ) Van Hulten-betänkandet är ett viktigt bidrag till arbetet i samband med reformeringen av EU och det arbete som genomförs av kommissionär Kinnock .
En effektiv och dynamisk kommission är en förutsättning för en utvidgad europeisk union .
Skyddet av EU : s ekonomiska intressen ingår som en del av dagordningen för reformeringen .
EPLP anser - samtidigt som vi håller med om att det finns behov av att förbättra skyddet av EU : s ekonomiska intressen - att förhållningssättet med tre steg för inrättandet av ett offentligt åklagarämbete på gemenskapsnivå , som beskrivs i betänkandet , inte är rätt sätt att gå vidare på och att det krävs en betydligt mer ingående diskussion för att hitta sätt att ta itu med bedrägeri som är effektiva i alla medlemsstater .
EPLP stöder endast inrättandet av ett offentligt åklagarämbete på gemenskapsnivå så som detta beskrivs i punkt 38 för att ge tillträde till information för att underlätta åtal - vid nationella domstolar - av de som gör sig skyldiga till bedrägeri med skattemedel .
EPLP anser också att ett inrättande av en kommitté om normer inom EU : s offentliga verksamhet skulle främja alla Europeiska unionens institutioner , inklusive Europaparlamentet .
( Sammanträdet avbröts kl .
13.20 och återupptogs kl .
15.00 . )
 
Fredsprocessen i Mellanöstern ( fortsättning ) Nästa punkt på föredragningslistan är fortsättningen på debatten om rådets och kommissionens uttalande om fredsprocessen i Mellanöstern . .
( EN ) Jag är mycket tacksam mot rådets ordförande för uttalandet i förmiddags om Mellanöstern i början av denna debatt och för en del av minister Gamas insikter , efter det han i största hast rest hit från regionen i fråga .
Det enda jag beklagar är att mitt initiativ till att öppna Europeiska återuppbyggnadsbyrån i måndags innebar att jag inte personligen kunde resa till Mellanöstern , även om , som jag nämnde tidigare - vilket är en annan historia - ödet såg till att strandsätta mig på Münchens flygplats i stället för att transportera mig till Thessaloniki .
Sånt är livet .
Jag hoppas att ledamöterna ursäktar om jag inte kan stanna hela debatten , vilket jag skulle ha gjort under normala förhållanden .
Debatten hade planerats till denna förmiddag och på grundval av detta hade jag arrangerat ett möte med besökare från Balkanområdet i kväll .
Jag hoppas alltså att kammaren visar förståelse i detta fall .
Jag kan försäkra er om att detta inte är något som jag kommer att göra till en vana .
I likhet med ledamöterna välkomnar jag Förenta staternas initiativ till att återuppta förhandlingarna mellan Syrien och Israel , trots syriernas beslut att det behövde mer tid innan de kunde återuppta samtalen som planerats att starta återigen i dag .
Det finns ett gott hopp om att det skall kunna gå att bygga en grund för ett fredsavtal inom den närmaste framtiden .
Jag hoppas också att framsteg i samband med förhandlingarna med syrierna kommer att bana väg för ett tidigt återupptagande av samtalen mellan libaneserna och israelerna , som sedan skulle kunna föras parallellt för att uppnå en övergripande överenskommelse rörande Israels förbindelser med dess grannländer i norr .
Samtidigt får vi inte glömma bort den palestinska sidan .
Palestiniernas situation har alltid utgjort själva grundfrågan i konflikten .
En rättvis och även storsint överenskommelse med dem är fortfarande nyckeln till en hållbar fred i Mellanöstern .
Israelerna och palestinierna har gjort betydande framsteg när det rör genomförandet av Sharm el Sheikhs samförståndsavtal .
Även om det skett en viss avmattning , antar jag att tillbakadragandet av de återstående israeliska trupperna snart kommer att ske .
På samma sätt , trots att tidtabellen för ramavtalet om permanent status i förgår förflyttades till en tidpunkt bortom tidsfristen i mitten på februari , hoppas jag innerligt att den mycket viktigare september-tidsfristen för det slutliga avtalet om permanent status kommer att uppfyllas .
Jag fick uppfattningen att detta också var premiärminister Baraks och ordförande Arafats ståndpunkt när de sammanträdde i måndags .
Ledamöterna skall veta att vi särskilt engagerar oss för att man skall återuppta de multilaterala samtalen om framsteg .
Detta är långt ifrån okomplicerat , men vi skall göra vad vi kan för att uppnå detta i nära samarbete med medarrangörer från Förenta staterna och Ryssland , såväl som med de regionala parterna .
Vi har ett särskilt ansvar för främjandet av den regionala ekonomiska utvecklingen .
Inledningen av samtalen med Syrien banade väg för ett sammankallande av den multilaterala styrgruppen i Moskva vid slutet av månaden .
Jag ser fram emot att få delta i detta sammanträde och hoppas att vi åtminstone kan börja se framåt igen .
Europeiska unionen har en viktig roll inom fredsprocessen , precis som alla sidor - palestinier , israeler , deras arabiska grannländer och Förenta staterna - har erkänt .
Vår roll är inte heller begränsad till att bara vara bank .
Vi måste vara beredda att handla snabbt för att stärka freden i regionen .
Men vi bör inte lura oss själva : Ett heltäckande fredsavtal i Mellanöstern kostar mycket i reda pengar .
Kommissionen håller redan på att bedöma konsekvenserna för Europeiska unionen av den senaste utvecklingen vad gäller främjande åtgärder .
Vi har för avsikt att snart meddela våra slutsatser i frågan till parlamentet och rådet .
Men låt mig påminna ledamöterna om att vi i Europeiska unionen inte är några slöfockar när det gäller ekonomiskt stöd till fredsprocessen .
Vi är den största biståndsgivaren av alla när det rör medel till palestinierna .
Vi har också erbjudit mycket omfattande stöd till Jordanien , Libanon , Syrien och Egypten .
Tillsammans med israelerna har vi upprättat ett närmare samarbete inom en rad områden som är av särskild betydelse för dem .
Gemenskapens bidrag på över 600 miljoner euro i stöd och lån mellan 1994 och 1998 , understödde den palestinska myndigheten på ett effektivt sätt och bidrog i hög grad till återuppbyggnaden av den förfallna fysiska infrastrukturen på Västbanken och i Gazaområdet .
Europeiska unionens medlemsstater bidrog tillsammans med ytterligare 860 miljoner under denna viktiga period .
Låt mig i detta sammanhang applådera de viktiga steg som den palestinska myndigheten nyligen vidtagit för förbättring av öppenheten rörande budgeten .
Ordförande Arafat kommer att sammanträda med ministerrådet nästa vecka .
Detta är ett bra tillfälle att ta itu med behovet av att vidta liknande djärva åtgärder för att förbättra den palestinska förvaltningen och stärka rättssäkerheten .
Kommissionen deltar aktivt i dessa ansträngningar .
Kommissionen har också ökat sitt planerade stöd till regionala samarbetsprojekt mellan israeler och araber .
Vi avsatte mer än 20 miljoner euro till sådana projekt under förra året .
Detta paket omfattade förnyat bistånd till mellanstatlig verksamhet och gränsöverskridande samarbete då israeler och araber träffas på icke-statlig och sakkunnignivå .
Ledamöterna känner till att Europeiska unionen är den största ekonomiska biståndsgivaren rörande övergripande initiativ för att uppnå en försoning mellan folken i Mellanöstern .
En rad frågor växer på ett naturligt sätt fram som ytterligare möjliga mål för stöd från gemenskapen under fredsprocessens kommande fas - bland dessa finns hjälp till att konsolidera en bosättning inom Golanområdet , både vad gäller bidrag till säkerhetsarrangemang och stöd till minröjning och återuppbyggnad av samhällen på Golanhöjderna .
Den syriska ekonomiska utvecklingen kommer att behöva stöd under övergången från en krigs- till en fredsekonomi .
Återuppbyggnaden och återanpassningen av södra Libanon , det enda området i Mellanöstern med en pågående militär konflikt , kommer också att kräva avsevärda ansträngningar .
Vi behöver också fortsätta att ge stöd till den ekonomiska reformeringen och den sociala utvecklingen i Libanon som helhet .
Det behövs en lösning på det palestinska flyktingproblemet - det är den största flyktinggruppen i världen och uppgår till nästan 5 miljoner personer - vilket visar litet av de enorma utmaningar som ligger framför oss .
Vi måste stödja initiativ som ökar tillgängligheten och förbättrar distributionen och förvaltningen av regionens mycket knappa vattenresurser .
Till sist det kanske mest viktiga - vi måste främja ett närmare regionalt samarbete inom en rad områden och föra samman alla berörda länder i ett gemensamt försök att ta itu med deras gemensamma problem .
Det är redan uppenbart att de ekonomiska resurser som för närvarande finns tillgängliga för bistånd till denna del av världen inte kommer att räcka till för det stöd som kommer att krävas i det fall man uppnår en permanent fred .
Jag vill betona detta .
Jag vill verkligen påminna rådet och , om det blir nödvändigt , parlamentet , att vi inte i fortsättningen bör tillåta att det uppstår en klyfta mellan vår retorik och vad vi faktiskt kan åstadkomma .
Jag upprepar att en förändring av Mellanösternpolitiken kommer att fordra en växling vad gäller det stöd vi kommer att tillfrågas om och förväntas tillhandahålla .
Låt mig tillägga att vi vill tillhandahålla detta .
Vi har nått framgångar under de senaste veckorna och månaderna , som minister Gama nämnde tidigare .
Men det kommer oundvikligen att bli en tuff process som kommer att innehålla svårigheter och besvikelser .
Vi kommer att göra allt som står i vår makt för att se till att processen slutar i framgång och för att följa de åtaganden och utmaningar som detta resultat leder fram till .
Låt mig slutligen upprepa för de som anlänt till kammaren under de senaste minuterna , vad jag sade i början : Jag kommer inte att kunna stanna till debattens slut , framför allt beroende på att jag hade antagit att debatten skulle ske i förmiddags och därför hade bestämt att delta i ett sammanträde om Balkanområdet i kväll .
Jag hoppas att kammaren kan visa förståelse för detta .
( Applåder ) ) Herr talman !
Vi förstår kommissionär Patten mycket väl .
Jag vill bara säga att förbindelserna med Madrid i vanliga fall är ganska så bra , och att jag därför snart hoppas få se honom där .
De uttalanden vi under dagens lopp har hört om fredsprocessen i Mellanöstern kommer mycket lägligt efter den pressande rundresa minister Gama - jag beklagar hans frånvaro - tillsammans med tre andra representanter från rådet gjorde i området .
De nyheter man rapporterat om i massmedia skulle kunna få oss att se pessimistiskt på situationen .
Jag tror ärligt talat att en utvärdering av det här slaget inte överensstämmer med verkligheten .
Jag delar därför kommissionär Pattens positiva inställning .
Jag skall förklara varför : Det är sant att den israeliska regeringen har flyttat fram det tredje överlämnandet till de palestinska myndigheterna av mark på Västbanken .
Men det är också sant att man sedan Sharm el-Sheikh har överlämnat 39 procent av Västbanken och två tredjedelar av Gazaremsan till Palestina och att - vilket är än viktigare - nämnda avtal fram till nu har följts till punkt och pricka , till och med uppskovet är ett prerogativ från den israeliska regeringens sida som förutsetts i Sharm el-Sheikh .
Förutsatt , givetvis , att det inte dröjer mer än tre veckor , vilket är vad premiärminister Barak har lovat .
Å andra sidan är beslutet att flytta fram den andra samtalsrundan , som inleddes i Shepherdstown av Arabrepubliken Syrien , tvivelsutan en viktig händelse , men jag är övertygad om att hoppet från den 3 januari inte kommer att gå förlorat .
Herr talman , det faktum att kammarens alla politiska grupper inställer sig till den här debatten , som alltid är kontroversiell , med ett resolutionsförslag som man enhälligt har bifallit tycker jag är avgörande för vår politiska vilja att bestämt stödja de pågående fredsförhandlingarna .
Med samma kraft tar vi avstånd från våldshandlingar för att lösa meningsskiljaktigheter , må vara djupa , parterna emellan .
Enligt min mening är detta en garanti för båda parter , såväl ur politisk som ekonomisk synpunkt , för de åtaganden som kan förväntas av Europeiska unionen när det gäller kostnaderna för den fred vi alla så hett eftertraktar .
För att kunna garantera säkerheten i området och för att kunna bidra till att mildra rådande sociala skillnader förnekar ingen att detta är absolut nödvändigt .
Men det uppmärksammar också Europeiska unionens krav på att politiskt få delta i processen , i enlighet med vårt ekonomiska stöd så att det offentliggörs på motsvarande sätt , eftersom inte heller vi gör anspråk på att vara bankirer .
Europaparlamentets ordförande och hennes kommande resa till området kommer tvivelsutan att bidra till detta .
Herr talman !
Jag vill tacka kommissionär Patten för en utförlig beskrivning .
Jag vill gärna säga att jag ansluter mig till den ton som Galeote Quecedo angav här .
Vi i parlamentet stöder starkt fredsprocessen i Mellanöstern .
Det är ju en fredsprocess som äntligen är på gång .
Trots svårigheter och förseningar , är det ändå en skillnad som mellan natt och dag om vi tänker på hur processen såg ut för ett år sedan .
Jag vill understryka fyra punkter .
För det första innehåller Sharm el-Sheikh-avtalet en konkret tidsplan som alla vet för genomförandet av Israels åtaganden ; det gäller då interimsavtalet samt Hebron- och Wye-avtalen .
Medan förhandlingarna om slutlig fredsuppgörelse har inletts , tror jag att det är viktigt att hålla isär de två .
Brist på framsteg i slutstatusförhandlingarna bör inte äventyra genomförandet av de tre ovannämnda interimsavtalen .
Vad vi behöver bevaka i detta sammanhang är hur det går med hamnen i Gaza , den nordliga transitrutten mellan Gaza och Västbanken , ytterligare frisläppande av säkerhetsfångar och genomföranden av de ekonomiska åtagandena .
Den andra punkten gäller Syrien .
Där är naturligtvis gränsfrågan central .
Hur förhandlingarna går där , vet vi inte ännu .
Det viktiga är emellertid att de har inletts .
En viktig fråga i sammanhanget är den framtida vattenfördelningen .
Golan svarar i nuläget för mellan en tredjedel och en sjättedel av Israels vattenförsörjning .
Den tredje aspekten är fredssamtalen i Syrien som är nära sammankopplade med frågan om israeliskt tillbakadragande från södra Libanon .
Enligt uppgift från UNIFIL , finns det nu konkreta tecken på att Israel förbereder ett tillbakadragande , vilket vi välkomnar .
Utestående tvistefrågor är naturligtvis även där vattenproblematiken och de libanesiska Palestinaflyktingarnas situation .
Min sista punkt gäller den kommande palestinska staten .
Den kan komma att utropas under detta år , med eller utan Israels stöd .
Regeringen Barak har låtit förstå att man är inställd på att sluta ett fredsavtal med en stat som motpart .
Även om inte förhandlingarna är avslutade i september detta år , finns det inga fördragsmässiga hinder mot att en palestinsk stat skall utropas efter detta datum .
I detta sammanhang är det då viktigt för oss som stöder tanken på detta , att det blir som kommissionär Patten sade , nämligen en stat med insyn och att det blir en demokratisk stat .
Det vill vi alla medverka till .
Herr talman !
Jag skulle gärna först och främst vilja hänvisa till den gemensamma resolution som skall läggas fram som avslutning på den här debatten och till vilken min grupp bidragit och som vi naturligtvis godkänner .
Mer specifikt vill jag dock uttrycka min glädje över att Israel och Syrien efter så lång tid återigen samtalar för att lösa sina meningsskiljaktigheter .
De nya förhandlingarna är i alla fall ett viktigt steg mot en varaktig fred i mellanöstern .
Därför är det synd att de här fredssamtalen skjutits upp tills vidare .
Båda parter kommer mycket riktigt att behöva göra stora insatser .
En varaktig fred i det här området kan förverkligas först genom ett avtal i vilket säkerheten för de israeliska gränserna och Syriens integritet kan garanteras .
För det behövs också fasta diplomatiska förbindelser och en oavbruten dialog .
Förutom de bilaterala mötena med Syrien hoppas jag att Israel inom överskådlig tid även skall inleda förhandlingar med Libanon och att en multilateral process skall visa sig möjlig inom ramen för det ekonomiska och regionala samarbetet .
Det är ändå beklagansvärt att Europeiska unionen , en av de viktigaste ekonomiska givarna , fortfarande inte kan spela en viktig politisk roll i fredsprocessen .
Den här fredsprocessen i Mellanöstern är en av prioriteterna för Europeiska unionens gemensamma utrikes- och säkerhetspolitik .
Här har Solana , den höga representanten i rådet , en särskild funktion .
Kommissionen och medlemsstaterna måste också uppmuntras att stödja projekt som kan hjälpa till att bygga upp förståelse och partnership mellan de olika folkgrupperna i det här området .
Jag måste också påpeka Barcelonaprocessens betydelse som ju måste ha ett positivt inflytande på det regionala samarbetet .
I det avseendet stöder vi Libyens deltagande , på villkor att landet erkänner de mänskliga rättigheterna , avstår från att ge stöd till terrorister och ger sitt fullständiga stöd till fredsprocessen .
Det kvarstår naturligtvis många olösta problem och obesvarade frågor , även med palestinierna .
Alla vet att fredsprocessen är en lång och tung process men vi är övertygade om att med nödvändig tillförsikt , med den oumbärliga politiska viljan och med den ihärdighet som behövs så kommer vi att nå vårt gemensamma mål , nämligen ett fredligt och välmående Mellanöstern .
Herr talman !
Det är glädjande att fredsförhandlingarna , trots vissa uppskov och problem , pågår såväl mellan Israel och Palestina som mellan Israel och Syrien .
Sanningens minut närmar sig .
Är Israel berett att följa FN : s resolutioner och återlämna de arabiska områden som erövrades 1967 i utbyte mot fred och säkerhet ?
Kommer Israel att låta palestinska flyktingar återvända eller få kompensation ?
Kommer Israel att dela med sig av Jerusalem och floden Jordans vatten ?
Kommer det fria Palestina att bli en fullt demokratisk stat och därmed pålitlig som fredspartner ?
Kommer Syrien att fullt ut acceptera Israels existens och införa demokrati och rättsstatlighet ?
Att huvudansvaret för fredsprocessen ligger på ockupanten Israel hindrar inte att också de arabiska parterna har ett stort medansvar .
Mellanösternfreden angår oss emellertid alla .
Därför är det bra att EU agerar som fadder till den palestinska staten .
Mot denna bakgrund vill jag avsluta med en märklig historia i EU-landet Sverige .
Där hålls en internationell regeringskonferens om Hitlers judeutrotning , vilket självklart är ett välkommet initiativ .
Bland fyrtiosju inbjudna stater från samtliga världsdelar finns emellertid inte en enda av de arabstater som ingår i EU : s Barcelonaprocess .
Detta har tolkats som att den arabiska hållningen gentemot Israel av européer skulle betraktas på samma sätt som nazismens antisemitism , vilket ju är fullständigt felaktigt .
Arabvärldens Israelkritik har byggt på samma sorts antikolonialism som exempelvis Algeriets frihetskamp mot Frankrike .
Men i dag har ju Egypten , Jordanien och Palestina fördragsfäst fred med Israel .
Därför undrar jag om inte kommissionär Patten håller med mig om att det hade varit rimligt och lämpligt att åtminstone någon arabstat hade varit inbjuden till förintelsekonferensen i Stockholm .
Herr talman !
Jag vill verkligen tacka kommissionär Patten för de kunskaper han gett prov på när det gäller svårigheterna i fredsprocessen och den utmaning som Europeiska unionen har antagit när det gäller att förverkliga den .
Det är verkligen dags för fred i Mellanöstern .
Det är dags att avsluta den epok i historien som inleddes med Balford-förklaringen 1917 och det arabisk-israeliska kriget 1948 .
Det är dags att det äntligen blir säkra gränser för samtliga länder i området , politiska , sociala och ekonomiska rättigheter , mänskliga rättigheter som erkänns och tillämpas i Syrien , Palestina och Israel , överallt .
Det handlar också om att varje folk och varje individ skall kunna leva självständigt och demokratiskt , men för att det skall kunna förverkligas är det nödvändigt att samtliga parter i konflikten har modet att tillämpa fred och rätt , att man erkänner den andre som en partner och inte som en undersåte som man måste bevilja eftergifter .
Jag tänker i första hand på knuten Palestina-Israel , men det gäller även de områden som ockuperades i Golan 1967 och den södra delen av Libanon efter 1982 .
Israel måste ta sitt ansvar , lämna de ockuperade områdena och dela på vattenresurserna , men samtidigt måste Israel få garantier för sin säkerhet och kunna leva i fred i ekonomiskt och politiskt utbyte med samtliga länder i området .
Men säkerheten gäller inte bara Israel .
Samma sak gäller de övriga länderna , i första hand palestinierna som fortfarande lever under militär ockupation och som fortfarande i dag , trots de avtal som undertecknats från och med Oslo , ser sin mark konfiskerad i områdena B och C. Efter Oslo och fram till och med den 17 oktober 1999 har 174 tusen dunans mark konfiskerats , varav 8 462 under den nya regeringen Barak .
Träd har ryckts upp med rötterna , hus har förstörts och framför allt i östra Jerusalem har utnyttjandet av vattnet inskränkts eller förvägrats , medan bosättningarna fortsätter och hela tiden ökar .
Det råder emellertid inget tvivel om att i och med att den nya regeringen valts så har framsteg gjorts , åtminstone har man börjat förhandla igen .
Men det kan inte finnas någon stabil och varaktig fred i Mellanöstern om inte palestinierna får sin egen stat , om de inte fritt kan röra sig på sitt eget territorium .
Det internationella samfundet måste helt enkelt tillämpa resolutionerna nr 332 , 248 , 245 och 194 .
Det är oroande att förbindelserna med Syrien har skjutits på framtiden , liksom Baraks beslut att skjuta upp tillbakadragandet av den israeliska armén och avtalen från Sharm el-Sheikh .
Det är utomordentligt viktigt att Europeiska unionen kan spela en politisk roll i förhandlingarna parallellt med sin roll när det gäller ekonomiskt bistånd .
Vi kan inte nöja oss med att stå i kulisserna , vi måste i stället spela en huvudroll , utan att för den skull hamna på kollisionskurs med USA , som minister Gama påpekade .
Herr talman !
Låt mig först uttrycka mina tack och min uppskattning till kommissionär Patten för hans kommentarer här i dag , särskilt i samband med Europeiska unionens roll i fredsprocessen och för att han bekräftar att vår roll inte bara innebär att vara " bank " för hela verksamheten .
Jag blev djupt besviken när jag fick höra nyheterna i veckan om att fredssamtalen mellan Israel och Syrien hade skjutits upp .
Jag hoppas verkligen att man kan nå en kompromiss , så att fredssamtalen snabbt kan återupptas .
Vi kan emellertid inte förneka att det skett en del positiva politiska framsteg i Mellanöstern under den senaste tiden .
Det faktum att den syriske utrikesministern och den israeliske premiärministern nyligen satt vid samma bord i Förenta staterna för första gången någonsin är ett tecken på går att övervinna det gamla hatet och fientligheterna .
De politiska ledarna måste visa verkligt mod för att anta en gemensam ram som kan leda fram till en övergripande fred i Mellanöstern .
Jag vet att om det går att nå ett avtal mellan Syrien och Israel , kommer Israels premiärminister att möta verkliga protester mot alla nya avtal med Syrien i framtida folkomröstningar .
Bosättarna på Golanhöjderna kommer att kräva kompensation och det måste bli garantier rörande säkerheten .
Om Syrien skulle vara redo att ta itu med säkerhetsfrågan , skulle utsikterna för en lösning på Israel-Syrienfrågan vara goda .
Vad gäller Palestinafrågan inser jag att det fortfarande finns vissa svårigheter rörande genomförandet av vissa aspekter av Wye-avtalet .
De största problemområdena omfattar för tillfället omstrukturering , såväl som överflyttning av territorier .
Den låga graden av frisläppande av palestinska fångar och det faktum att den israeliska regeringen verkar stoppa tillämpningen av byggnadstillstånd som redan beviljats , såväl som att inte utfärda nya , utgör ytterligare hinder .
Dessa frågor har uppenbarligen hejdat framstegen i förhandlingarna om den permanenta statusen , även om - tror jag - dessa samtal inte kommer att stoppas för evigt .
Den största svårigheten just nu när det gäller att få igång förhandlingarna , verkar vara att palestinierna vill att man först och främst skall lösa gränsfrågan , medan den israeliska regeringen säger att denna endast kan lösas om man först når en lösning i frågan om bosättningarna och säkerheten .
För tillfället verkar det som om båda sidor har accepterat att man inte kan komma överens om någonting , förrän man kommit överens om allt .
Medan , sammanfattningsvis , andra länder i Mellanöstern haft betänkligheter rörande fredsprocessens allmänna riktning , nu när den syriska regeringen också deltar i fredsprocessen , är Egypten och andra länder i regionen redo att gå vidare .
Jag hoppas verkligen att - när det gäller att förbättra säkerheten och livskvaliteten för folken i Mellanöstern - alla tongivande parter så snart som möjligt ser till att ingå ett övergripande avtal om alla viktiga frågor som behöver få en lösning .
Herr talman , ärade kolleger !
De olika resolutionsförslag som lagts fram i parlamentet ger en god bild av läget i Mellanöstern .
Det finns de som applåderar nya avtal mellan Israel och Syrien , men bara någon enstaka riktar uppmärksamheten mot det verkliga och centrala problemet när det gäller Mellanöstern .
Ögonblicket är nu inne , ärade kolleger , att lösa upp en av knutpunkterna när det gäller den globala jämvikten .
Ögonblicket är nu inne för Israel att hålla sina gamla löften och slutgiltigt dra sig tillbaka från de områden man ockuperat och slutgiltigt och en gång för alla erkänna den palestinska myndigheten , vars återupptagna diplomatiska verksamhet utan tvekan kommer att ha en framtid så länge den befinner sig i Yasser Arafats erfarna händer .
Det är lika viktigt att vi inte förlorar den irakiska frågan ur sikte , en fråga som ingen längre talar om utan man förtränger problemen för miljontals kvinnor , gamla och barn , offer för ett embargo som är lika arrogant som gement .
Jag vet inte vad Syrien och Israel verkligen skulle vilja eller skulle kunna göra , men jag vet att vår institution skulle kunna göra mycket och det är på tiden att vi ägnar oss åt hur människor lever med samma kraft vi som vi ägnar oss åt tändanordningarna till våra lika kalla som vaga och artificiella neonlampor , som kan lysa upp ett hus , men verkligen inte världen under tredje millenniet .
Herr talman !
Den israeliska författaren , Amos Oz , beskrev nyligen mycket träffande det kyliga förhandlingsklimatet mellan Israel och Syrien .
Oz hade fått intrycket att syrierna ansåg att de i utbyte för Golanhöjden endast behövde faxa ett mottagningsbevis till israelerna .
Den tanken av Oz dyker också upp i den israeliska pressen .
Den återger kontrasten mellan premiärminister Baraks personliga fredsansträngningar och den reserverade hållningen , den rent av fysiska frånvaron , hos Damaskus starke man , president Assad , vid förhandlingsbordet i Förenta staterna .
Det var väl ändå Assad som skulle vara Baraks samtalspartner och inte hans utrikesminister .
När det gäller minister Farouk al-Sharas beteende i Shepherdstown är israelerna mycket upprörda .
Hans hållning gentemot premiärminister Ehud Barak var rent ut förnedrande .
Vadan denna uppmärksamhet för elementära diplomatiska umgängesformer i en seg territoriell förhandlingsprocess ?
Jo , syrierna förstör bara för sig själva .
När allt kommer omkring är det de israeliska väljarna som skall uttala sig om huruvida Golanhöjderna skall lämnas tillbaka .
I alla resolutioner som lagts fram uttalas en djup önskan om en större europeisk roll i fredsprocessen .
Det är dock frågan om Bryssel kan skaffa fram de miljarder dollar som de israeliska och syriska myndigheterna är ute efter hos sin fredsbeskyddare , Förenta staterna .
Då talar vi ändå inte om de tunga , lika dyra säkerhetsgarantierna om Israel drar sig tillbaka från Golan .
Slutligen en fråga till rådet och kommissionen .
Vad är sant i pressens uppgifter om att det portugisiska ordförandeskapet redan utlovat trupper till en fredsbevarande styrka i Golan ?
Herr talman !
Sanningen är att brytningen eller förseningen sine die av de pågående samtalen mellan syrier och israeler inte är en bra nyhet .
Det är inte heller en bra nyhet att ett nytt bombattentat inträffade i förrgår och 16 personer skadades .
Det är tydligt att Förenta nationerna för en gång skull inte har lyckats i sina medlingsförsök , och det är faktiskt svårlösta hinder .
Syrierna försöker än en gång att få Golan under sin suveränitet och jurisdiktion och få tillbaks de gränser som gällde före den 4 juni 1967 medan israelerna vill ha gränserna dragna som de var 1923 , eftersom det är bättre för dem .
Avbrottet i samtalet mellan syrierna och israelerna är inte den enda förseningen i fredsprocessen i Mellanöstern .
Just nu har tillämpningen av ramavtalet mellan Palestina och Israel också hävts .
Efter samtalen i förrgår mellan Israels premiärminister och Palestinas ledare begärde den israeliska premiärministern en två månader lång ajournering från och med den 13 februari , sista dag för verkställandet av ramavtalet om situationen på Västbanken och Gazaremsan .
Vad kan Europeiska unionen göra i en sådan här situation ?
Inte mycket , tyvärr .
Vi måste givetvis stödja förhandlingarna ledda av Förenta staterna .
Vi måste intensifiera våra kontakter .
Europeiska unionens sändebud , ambassadör Moratinos , har inom ramen för Europeiska unionens befogenheter utfört sitt uppdrag med stor omsorg och effektivitet .
Detta till trots kan vi ana en viss maktlöshet , när de båda förhandlingspartnerna i helgen tar flyget hem till Förenta staterna får vi inte förglömma att för varje 100 dollar som spenderas i fredsprocessen kommer 60 från Europeiska unionen .
När vi dessutom beaktar att nästa möte kommer att hållas i Moskva , så blir Europeiska unionens närvaro något patetisk .
Inför det portugisiska ordförandeskapet insisterar jag på en mera central roll , det är dags för Europeiska unionen att ta över och bli mera delaktig .
Jag hoppas att nästa besök i regionen av Europaparlamentets talman , samt av de interparlamentariska delegationerna och deras ordförande , tillåter oss att inleda en mera initiativrik etapp där Europeiska unionen tydligare kan delta i denna komplicerade och svåra fredsprocess .
Herr talman , herr rådsordförande , kommissionär Patten !
Jag vill tacka för era redogörelser , särskilt gäller det kommissionär Patten vars analys jag helt och fullt delar .
Jag kommer av den anledningen ej att upprepa något av vad han sagt .
I stället vill jag göra tre kommentarer som kommissionär Patten måhända har samma syn på men som han av olika skäl inte kan formulera lika öppet som en ledamot kan göra .
Det första är att jag tror att vi har anledning att glädja oss över det avtal som finns mellan Israel och den palestinska myndigheten för självbestämmande .
Nu finns det dock tillräckligt med avtal : Oslo , Wye Plantation , Sharm-el-Sheik .
Det räcker så , nu måste de uppfyllas också .
På den punkten delar jag emellertid min kollega Salafrancas skepsis när han säger att det kom dåliga nyheter från Israel , närmare bestämt att även detta senaste avtal inte kommer att kunna uppfyllas i tid .
Den andra punkten gäller återupptagandet av förhandlingarna mellan Syrien och Israel .
Detta är , menar jag , en högst glädjande nyhet .
Men denna vecka har vi också fått höra att Barak inte reser till Washington och att förhandlingarna därmed inte kan fortsättas .
Jag vill klart och tydligt slå fast att om Golanhöjderna lämnas tillbaka till Syrien så är problemet löst i denna region .
Gällande frågan om folkomröstning som berörts av flera kolleger : Vi måste nu fråga oss om man verkligen alltid måste hålla folkomröstning för att kunna uppfylla förpliktelser ur internationell rätt och folkrätten .
I Tyskland skulle man förmodligen glädja sig mycket om vi sade att vi genomför en folkomröstning för betalningen till Europeiska unionen ; men vi gör det oberoende av huruvida det tyska folket är villigt att betala .
Det skulle vara en likartad situation .
Min tredje och sista punkt gäller Europeiska unionens roll .
Här vill jag verkligen framhålla den enastående roll som det särskilda sändebudet Moratinos har spelat i regionen , samt även det vi åstadkommit i form av finansiering , kommissionär Patten .
Ni skall veta att ni alltid kan få stöd för ert förslag i detta parlament .
Vi kommer att finnas där när det skall finansieras .
Vi bör dock också spela en politisk roll , som ju Moratinos inte kan göra helt själv i denna region .
Rådsordförandeskapet måste då aktiveras , Mister GASP måste då ta sig till regionen , och vi måste själva bjuda in förespråkarna för fredsprocessen , på samma sätt som ryssarna gjort .
Då har vi tagit det ansvar som motsvarar vårt engagemang och bidrag .
Herr talman , kommissionär Patten , kära kolleger !
De senaste fredsförhandlingarna som inletts i Förenta staterna mellan Israel och Syrien är en vändpunkt i Mellanösterns historia , en vändpunkt som man väntat på i femtio år nu och som uppenbarligen är svår att förhandla om .
Det blir inget möte i dag i Shepherdstown , men vi skall hoppas , såsom kommissionär Patten nyss sade , att detta uppskjutande av förhandlingarna på grund av de senaste kraven från Syrien , bara är en incident på vägen mot ett fredsavtal som kan ändra hela Mellanösterns utseende .
Det är vad vår resolution uttrycker : en förhoppning om ett rimligt och rättvist avtal , grundat på respekt för de suveräna staterna och rätten att leva i säkerhet inom säkra och erkända gränser .
Alla utländska trupper , inbegripet de syriska , måste alltså lämna Libanon , i enlighet med resolution 520 från Förenta nationernas säkerhetsråd .
Kan vi hoppas på att vi i juli 2000 - det datum som Ehud Barak lovat - fått uppleva en israelisk reträtt ur södra Libanon ?
Kan unionen hoppas på ett dubbelt fredsavtal mellan Israel och dess grannar i norr ?
Vi tror det .
Vi vill tro det .
Aldrig har parternas beslutsamhet varit starkare .
Jag skulle också vilja betona en punkt som förefaller mig grundläggande : balansen som måste känneteckna vårt europeiska budskap , en politisk balans mellan dem som deltar i förhandlingarna naturligtvis , men också balans mellan befolkningarna .
Efter attentatet mot Hadera i måndags måste vi upprepa vårt fördömande av varje form av terrorism .
Och apropå balans , eller obalans snarare i detta sammanhang , skulle jag vilja lägga till hur beklagligt det är att återigen tvingas konstatera vilken svag politisk roll Europa spelar när det gäller att lösa konflikten .
Vid lunchtid i dag tog rådets ordförande Gama upp Europas ekonomiska och handelsmässiga stöd till regionen .
Man måste trots allt konstatera att inledandet av fredsprocessen för närvarande i huvudsak är Washingtons verk .
Syrierna har , liksom andra arabiska länder före dem , valt ut amerikanerna för att beskydda förhandlingarna .
Det är också det val den hebreiska staten gjort där Europa , det är ett faktum och inte någon bedömning , lider av en partisk offentlig bild .
Det är alltså rätt tillfälle att på nytt säga till kommissionär Patten , till Solana och till Moratinos , att vi verkligen räknar med deras ansträngningar för att den europeiska rösten skall höras , i strävan efter en fredlig lösning av konflikten .
Och även om det är svårt för Europa att tala med en röst om fredsprocessen kan , och måste vi , ändå tala om den i samma anda av förtroende och solidaritet .
Herr talman !
Jag tror att det i denna fråga finns , trots de olika nyanserna , en allmänt samstämmig syn i Europaparlamentet , liksom jag också tror att de flesta instämmer i de allmänt positiva ståndpunkter som Patten redogjorde för .
På de få sekunder som står till mitt förfogande skulle jag vilja understryka en punkt som nästan alla talare har tagit upp , det vill säga frågan om Europas nedgraderade och politiskt svaga roll .
Kravet på att uppgradera Europas roll har inte framförts bara för att även vi skall spela en roll och delta , för att få ta del av Förenta staternas glans , utan på grund av , tror jag , att det finns en patologi mot den amerikanska politiken , som beror både på den enögdhet med vilken landet betraktar många frågor i Mellanöstern och på dess relation till de olika länderna , som Irak , Libyen , Syrien , men även på att landet bedriver en politik som tar liten hänsyn till de grundläggande principerna i den internationella rätten .
Europeiska unionen skulle kunna bedriva en politik som var mycket mer konkret , energisk och dynamisk och som grundade sig på de beslut som hittills har fattats av FN .
I den meningen tror jag att vissa punkter , som till exempel frågan om Israels tillbakadragande från de områden som landet erövrade 1967 , är nyckelpunkter på vilka Europa skulle kunna spela en roll och frigöra en mer allmän och positiv dynamik .
Herr talman , herr kommissionär , ärade damer och herrar !
Den israeliska fredsprocessen har gått i baklås innan den ens kommit igång på allvar .
Tyvärr !
Detta är dock inte särskilt överraskande och inte heller något att oroa sig över ; men det visar vikten av att Europeiska unionen och även Europaparlamentet stöder den fredsprocess mellan Israel och Syrien som lamslogs för fyra år sedan och som utgör en av grundförutsättningarna för fred i Mellanöstern .
Med tanke på den säkerhetspolitiska dimensionen i fredsprocessen är tålamod på sin plats .
Att president Clinton gärna skulle se en utrikespolitisk framgång i Mellanöstern mot slutet av sitt tjänstetid är begripligt , men får förstås inte leda till ett överilat förhandlingsresultat .
Om Europeiska unionen skall räknas som den största bidragsgivaren i regionen och vill tas på allvar i politiken krävs inte bara att man talar med en enda röst utan framför allt en viss balans .
Europeiska unionen måste undvika att bli betraktad som partisk .
Något som man inte alltid lyckats med i det förflutna .
Av den anledningen är man inte heller i någon högre grad tongivande i Mellanöstern .
I detta sammanhang måste jag ställa frågan hur samordnad Europeiska unionens utrikespolitik i själva verket är .
Denna fråga infinner sig inte bara i samband med rolluppdelningen mellan kommissionens kommissionär för utrikespolitik Chris Patten och Mister GASP Javier Solana , utan även med tanke på kommissionens ordförande Prodis inbjudan till Libyens statschef Khadaffi .
Jag erinrar mig den i Mellanöstern utomordentligt aktive före detta österrikiske förbundskanslern Kreisky ; genom att bjuda in Khadaffi orsakade han på sin tid för många år sedan mer skada än nytta .
När det gäller den säkerhetspolitiska dimensionen av återlämnandet av Golanhöjderna måste EU göra klart att ett sådant steg måste komma mot slutet av fredsprocessen med Syrien och inte i början .
Syriens motprestation får dock inte inskränka sig till en normalisering av de diplomatiska förbindelserna till Israel .
Till och med i en tidsålder då raketer når överallt måste faran att israeliskt territorium kan bli beskjutet från Golanhöjderna så som skedde 1967 avvärjas .
För detta ändamål krävs ett effektivt övervakningssystem .
För det andra måste en fred med Syrien i slutändan också leda till fred med Libanon .
Den israeliske ministerpresidenten Baraks uppställda mål att dra tillbaka de israeliska trupperna från säkerhetszonen i södra Libanon till juli år 2000 måste understödjas .
Emellertid måste också Syrien vidta motsvarande åtgärder ; landet har fortfarande en betydande truppnärvaro i Bekaa-slätten i Libanon och utövar även ett inflytande på terrororganisationer i Libanon .
Det åligger Syrien att strypa åtminstone delar av terrorscenen i Libanon .
Att detta kräver brådskande åtgärder visas av det senaste terrordådet i norra Israel .
Tidpunkten för en fred mellan Israel och Syrien är gynnsam , för även statschef Assad lär med tanke på sin ålder vilja lämna över ordnade förhållanden till sin efterföljare , läs sonen .
Därtill fattas en grundförutsättning , nämligen en demokratisk grundläggande ordning .
I stället kan EU erbjuda sin modell att genom ekonomisk-politisk sammanflätning , öppna gränser och frihet från tullbarriärer åstadkomma fred ; det är en modell som måste framställas som attraktiv över hela Mellanöstern .
Herr talman , herr kommissionär !
Vi är i denna debatt och i denna resolution medvetna om att det fortfarande återstår många hinder på vägen mot ett fullständigt förverkligande av fredsprocessen i Mellanöstern .
Men vi litar ändå på att den fredsvilja som folken i regionen visat kommer att segra och vi uppmanar Europeiska unionen att bidra genom att på nytt engagera sig .
Vi vill erinra om att unionen har spelat en roll i sammanhanget - vi har påmints om ambassadör Moratinos arbete , besöket av det portugisiska ordförandeskapet och nästa möte i Moskva - men vi skulle önska att det var kraftfullare .
Även om det har tillkommit nya problem under de senaste dagarna öppnar de återupptagna förhandlingarna mellan Syrien och Israel nya positiva framtidsutsikter och det är nödvändigt att handlingar följer på de beslut som fattades i Sharm el-Sheikh .
I vår gemensamma resolution erinrar vi om att de olösta frågor som återstår fortfarande är många och komplexa , kanske de mest komplexa - detta har mina kolleger redan påmint om - och till detta skall läggas det faktum att Libanon fortfarande inte sitter med vid förhandlingsbordet .
Europeiska unionen borde med andra ord ställa sig vid USA : s sida som en aktiv part i förhandlingarna och göra en kraftfull politisk satsning som tar fasta på framtiden för hela Medelhavsområdet och regionens oupplösliga band med Europa .
Unionen måste ingripa , eftersom instabilitet , krig och fattigdom i området redan har fått återverkningar på oss och får en allt större betydelse för vårt eget politiska , ekonomiska och sociala projekt .
Jag hoppas också att kommissionen och rådet skall agera mer samstämmigt och att Medelhavsområdet i dag blir ett högprioriterat område för Europeiska unionen .
Om man gör en ärlig analys av utvecklingen av Barcelonaprocessen så måste man erkänna att Europas uppmärksamhet i fråga om utvidgningen riskerar att delegera politiken i det området till den byråkratiska vardagslunken i pågående program och gällande bilaterala avtal .
Men framstegen i fredsprocessen , den politiska utvecklingen i många av de länderna , samt försöken att återuppliva de regionala organisationerna , som till exempel den arabiska Maghrebunionen , antyder att tiden kan vara inne för en ny dynamik i partnerskapet Europa-Medelhavet .
Kraftigt förenklat , kära vänner i rådet och kommissionen , är det budskap som vi vill skicka er att trots de ekonomiska åtagandena , som är viktiga , så är EU : s politiska roll fortfarande inte i nivå med den utveckling som pågår och som kan skönjas , såväl i Mellanöstern som i hela Medelhavsområdet .
Herr talman , kära kolleger !
Jag skulle i min tur vilja börja mitt personliga inlägg med att också jag gläds åt att Israel på nytt inlett fredsprocessen med palestinierna och syrierna .
Det är det påtagliga beviset för den oförsonliga viljan hos Ehud Barak och hans regering , att skapa fred under säkerhet .
Vi vet alla att ingenting någonsin är enkelt , och vi skall inte ta ut segern i förväg .
Oavsett förhandlingsläget är allt fortfarande möjligt , såväl det bästa som det värsta .
Det är anledningen till att jag , när det gäller Europa , personligen skulle vilja föreslå tre saker : till att börja med att vi européer försöker sluta upp med att hela tiden tjata , som vi säger på franska , vara smakdomare eller dela ut bra eller dåliga poäng .
Jag skulle vidare vilja att vi inte längre alltför mycket använder oss av korta turnéer i Mellanöstern , för övrigt ofta i Madeleine Albrights kölvatten .
Jag skulle framför allt också vilja att vi inleder en fördjupad diskussion med alla parter , och särskilt med israelerna , för att noga bedöma deras förhandlingsutrymme och fastställa de exakta punkter som vi kan trycka på .
För detta måste vi personligen träffa Ehud Barak , eftersom han är den som har nyckeln till freden i sin hand .
Och jag är säker på att våra vänner palestinierna sannolikt skulle föredra ett Europa som är mer förstående gentemot Israel , men som samtidigt , på samma sätt som Förenta staterna , skulle kunna utöva press för att avhjälpa vissa situationer .
Herr talman !
Jag avslutar med att säga att det är dags att sluta upp med att beklaga sig över vår svaga politiska styrka .
Om vi vill övergå från observatörsstatus till att bli aktörer måste vi vara beredda att betala det politiska priset för det .
Herr talman !
Jag vänder mig speciellt till det portugisiska ordförandeskapet och välkomnar Portugal som nytt ordförandeland för Europeiska unionens ministerråd .
Jag tror att Europas roll i Mellanöstern i framtiden kan finna en ny väg .
Europa måste på samma sätt som USA kunna vara trovärdigt , vinna respekt och få ett brett folkligt stöd bland medborgare och väljare i Mellanösterns enda demokrati - Israel .
Vi har ett förtroendekapital att bygga upp bland Israels medborgare .
Vi kan se på ett land som står utanför EU , t.ex.
Norge , som genom statsminister Kjell Magne Bondevik och utrikesminister Knut Vollebaek på ett förtroendeskapande sätt fortsatt att ha goda relationer med både Israel och med den arabiska sidan .
Man har det inte bara med Israels regering , utan även med Israels folk .
Vi kan också lära av Nederländerna och deras vattenprojekt .
Jag tror att Portugal som ordförandeland i EU har allt att vinna på att i EU : s namn jobba med vattenförsörjningsfrågorna som en av EU : s absolut centrala uppgifter i Mellanöstern .
Låt mig avsluta med att säga följande : Israel är Mellanösterns enda demokrati .
Låt oss aldrig glömma i vår kamp för demokrati , politisk pluralism och mänskliga rättigheter att Israel är en förebild och att Syrien med Hafez el-Assad är en av regionens absolut värsta diktaturer .
Herr talman !
Precis som det sägs i resolutionen om den överenskommelse som nåtts i den fråga som sysselsätter de flesta av kammarens grupper , så måste Europeiska unionens finansiella åtaganden i Mellanöstern åtföljas av en klar och tydlig politisk närvaro och unionen måste få delta i alla fredsförhandlingar .
Under årtionden - nästan så länge som stridigheterna har varat - har stora delar av allmänheten i Europa mobiliserat sig för att stävja hat och oförnuft och få det att ge vika för klokhet , enighet och sunt förnuft parterna emellan .
Folkets vilja har emellertid inte haft någon proportionell återverkan på de europeiska institutionerna .
Nämnvärda uttalanden i frågan har gjorts , som exempelvis Venecias , men de har fört en tynande tillvaro under årens lopp .
Denna politiska frånvaro , bristen på en verklig politisk vilja att agera samtidigt som det finns alltför många nationella röster av en annan mening , skadar inte bara unionen i det gemensamma europeiska projektet utan många utomeuropéer känner sig svikna , man skulle gärna se att vi tog på oss ett större ansvar och fick bättre samordning mellan utrikespolitik och annan politik .
Jag frågar såväl mig själv som er , ärade företrädare från rådet och kommissionen , om den nyligen inrättade tjänsten som GUSP : s höge representant kommer att åtföljas av en verklig enhetlig och gemensam politisk vilja .
Herr talman !
Europa kan inte påstå att det drar upp politiska framtidsutsikter i Mellanöstern och samtidigt blunda för viss verklighet , även om den är obehaglig .
Den första januari 2000 krävde Iran att staten Israel skulle upplösas , precis som Khadaffi , som Prodi ändå planerar att träffa inom kort , vilket skulle vara ett misstag .
Och när jag läser : upplösning av den judiska staten hör jag ekot av utrotning av det judiska folket .
Vi önskar alla av hela vårt hjärta att freden skall konkretiseras tillsammans med Iran , och absolut inte emot eller utan detta stora land .
Jag erinrar emellertid om att mellan Europa och Iran finns ändå dessa 13 fängslade judar som vi i stort sett inte vet någonting om , förutom att de riskerar döden .
Vi har tagit initiativ till förmån för dem , och vi kommer att ta ytterligare initiativ .
Vi kan slutligen inte fortsätta att låta bli att reagera när vi i pressen läser att de europeiska allmänna medlen skulle användas inom palestinskt territorium på ett minst sagt olagligt sätt , som de inte alls var avsedda för .
Det är kring den ekonomiska och kulturella utvecklingen som freden skall byggas .
Det är endast till detta som gemenskapens medel skall användas och jag kräver att kommissionen inleder en utvärdering som man sedan visar upp för parlamentet inom sex månader .
Jag har i enlighet med artikel 37.2 i arbetsordningen mottagit sex resolutionsförslag .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon .
 
Området frihet , säkerhet och rättvisa Nästa punkt på föredragningslistan är muntliga frågor till rådet ( B5-0040 / 99 ) och till kommissionen ( B5-0041 / 99 ) från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor om årsrapporten 1999 och om området frihet , säkerhet och rättvisa ( artikel 39 i Maastrichtfördraget ) .
Herr talman ! 1999 var det år då Amsterdamfördraget trädde i kraft , då Schengenavtalet införlivades och det extraordinära rådsmötet i Tammerfors hölls .
Det var här som rådets politiska vilja att inrätta området frihet , säkerhet och rättvisa inom Europeiska unionen som bäst kom till uttryck .
Rådet har beslutat sig för att utforma ett dokument för medborgarnas mänskliga rättigheter , vilket vi är glada över .
Man har beslutat sig för att införliva artikel 13 i fördraget , kampen mot all form av diskriminering och främlingsfientlighet , och man har beslutat sig för att harmonisera lagstiftningen om villkoren för mottagande och uppehållstillstånd samt garantera invandrarna en rättvis behandling likvärdig den som ges unionens övriga medborgare .
En politisk överenskommelse har också slutits - vilket vi tackar för - för de första förslagen om civilt samarbete .
Det här året har de rättsliga frågorna och inrikesfrågorna givits en politisk gemenskapsram .
Uppdraget har fallit på en och samme kommissionär , Antonio Vitorino , vilket vi tackar för .
Han har dessutom fått i uppdrag att konstruera en kontrollapparat för att mäta de reella framsteg gemenskapen har gjort inom det här området , men även medlemsländernas framsteg , vilket jag tycker är viktigt .
Vi tackar rådet för de här besluten , trots att Amsterdamfördraget för oss i kammaren innebar en viss besvikelse , det vill säga beslutet att låta vår roll anstå med fem år , vår möjlighet att aktivt delta , att demokratiskt kontrollera området frihet , säkerhet och rättvisa , liksom EG-domstolens roll i det hela .
Om vi tittar på de framsteg som gjorts under 1999 , vilket enligt fördraget åligger parlamentet , måste vi lämna de stora uttalandena och gå in på redan tagna och genomförda beslut och , herr talman , då mörknar panoramat rejält .
Det är som om rådet hade mer än ett ansikte och två händer , det som den ena undertecknar och uttalar sig om förkastar den andra .
Trots alla åtaganden på högsta nivå har rådet inte lyckats fatta de beslut man hade föresatt sig .
Programmen blir allt fler och de lappar över varandra och det finns ingen möjlighet att kontrollera genomförande- och effektivitetsnivån , parlamentet klara i alla fall inte av det .
Vi har vidarebefordrat ett antal frågor till rådet och jag vet att det är det portugisiska ordförandeskapets vilja att besvara var och en av dem .
Jag hoppas att rådet ändrar sin inställning till oss i kammaren från och med det här ordförandeskapet .
Det finns ingen egentlig överensstämmelse mellan rådets beslut och den politik som bedrivs .
Min grupp tvivlar , och kammaren tvivlar , på något som borde vara en god nyhet : införlivandet av Schengen i gemenskapsramen .
Schengen har , som vi tidigare nämnde , rigoröst införlivats , men på ett föga genomblickbart sätt .
Ingen information , inte en enda fråga har hamnat hos Europaparlamentet under förfarandets gång , varken om associeringen med Förenade kungariket eller Greklands införlivande eller förhandlingarna med Norge och Island .
Sak samma när det gäller immigrationspolitiken .
Vi har tillbringat vår tid med att utarbeta en mängd betänkanden , men vi vet inte vad som har hänt med initiativen .
De har försvunnit .
Vi får hoppas att år 2000 blir det år när allt genomförs , precis som 1999 var förväntningarnas år .
Vi får också hoppas att rådet gör en kraftansträngning och underställer sig kammarens kontroll .
Rådet har beslutat att rättsliga frågor och medborgarrätt skall vara en del av unionen .
Rådet kan agera i enlighet med sina beslut eller fortsätta att ömkligt vingklippa övriga institutioners delaktighet i detta betydelsefulla projekt .
Väljer man det sistnämnda bör man veta att det medför risker och kan komma att försvaga den grund området frihet , säkerhet och rättvisa vilar på .
Jag tror att vi i stället skulle kunna acceptera erbjudandet om ett avtal mellan institutionerna , så att vi kan gå vidare på ett annat sätt .
Fullgör med råge era skyldigheter gentemot parlamentet och förbered på det sättet framtiden .
Förse Europeiska kommissionen med erforderliga medel och det erkännande som behövs för att man skall kunna göra sitt arbete och för att man skall kunna kontrollera de framsteg som görs inom gemenskapen och i medlemsländerna .
Då får vi ett råd som håller måttet enligt de beslut som togs i Tammerfors för att få en friare , säkrare och mera rättvis union .
( Applåder ) , rådet .
( PT ) Herr talman , ärade ledamöter , herr kommissionär !
Det är med en viss sinnesrörelse jag nu i egenskap av medlem i rådet återvänder till detta parlament .
( Applåder ) Jag var en av de första portugisiska ledamöterna som 1986 tog de första stegen i den portugisiska integrationen i Europeiska unionen , och jag måste säga er , ärade ledamöter , herr ordförande , att den erfarenhet jag fick här , den politiska erfarenheten , var oerhört viktig i mitt liv , och den informationen och det bidrag vi alla kunde ge till det europeiska bygget präglade på ett avgörande sätt de år som jag tillbringade här , de präglade definitivt mitt liv .
Det är därför med stolthet och tillfredsställelse som jag befinner mig här , då jag har kunnat återse några av kollegerna från den tiden som fortfarande är kvar här i parlamentet .
Detta för att säga att det portugisiska ordförandeskapet - och jag själv och justitieministern , ansvariga för det rättsliga området - tillsammans med detta parlament vill inleda en ny period , främja en förbindelse mellan rådet och parlamentet vilken kommer att präglas av min parlamentariska erfarenhet i Europaparlamentet och givetvis också av de nationella parlamentariska erfarenheter som den betydelsefulla ledamoten i det nationella parlamentet fram till nu , justitieministern och min kollega har .
Ett första steg togs när vi träffades innan det portugisiska ordförandeskapet hade inletts , med ordföranden och vice ordföranden i utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor i Bryssel .
Vi fick möjlighet att bjuda in utskottets ordförande , ledamoten Watson och några av utskottsmedlemmarna till Lissabon , och vi redogjorde för våra synpunkter angående det portugisiska ordförandeskapets arbete på detta område .
Vi gjorde då vissa åtaganden som jag här mer formellt vill upprepa : Under alla möten med utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor , kommer en politisk företrädare för rådet , alltså inte en tjänsteman utan en företrädare för rådet på politisk nivå , någon från vår ministär , att hela tiden följa utskottets arbete ...
( Applåder ) och varje gång utskottet önskar det och på begäran av ordföranden , kommer jag själv och min kollega justitieministern att komma till Bryssel för att delta i mötena .
Redan i dag kommer vi att ge ordföranden för utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor den preliminära dagordningen för rådsmötet i mars och i maj , så att det i förväg kan sätta sig in de ämnen som kommer att diskuteras .
När det gäller 1999 , här har vi den speciella situationen att göra en utvärdering av det tyska och det finländska ordförandeskapet , skulle jag kunna börja med att säga att , utan att det inverkar på det skriftliga svar som i slutet av dessa arbeten kommer att överlämnas till ledamoten Ana Terrón i Cusí , som här lade in en protest för utskottets räkning , oberoende av de svar vi ger här , kommer ledamoten att få ett skriftligt svar .
Oberoende av detta skulle jag vilja säga att 1999 var ett betydelsefullt år i rådets arbete med de rättsliga och inrikes frågorna .
Samarbetet i de rättsliga och inrikes frågorna präglades av de långtgående förändringarna som genomfördes i Amsterdamfördraget och givetvis av införlivandet av Schengenavtalet i unionen .
Det tyska ordförandeskapet , vi måste erkänna detta , och säga det , hade en viktig roll i övergången från Maastrichtsystemet till Amsterdamsystemet .
Därefter kom starten för Europol-verksamheten i början av det finländska ordförandeskapet 1 juli 1999 .
Sedan hade vi en tredje viktig aspekt : toppmötet i Tammerfors , ett Europeiska rådet som helt ägnade sig åt rättsliga och inrikes frågor .
Toppmötet i Tammerfors präglades av en ny anda och av viljan att sätta området med frihet , säkerhet och rättvisa högst upp på den politiska dagordningen med ett bejakande av att den bör ligga kvar där .
Det som det portugisiska ordförandeskapet här återigen säger är att frågorna i samband med området med frihet , säkerhet och rättvisa genom vår vilja kommer att befinna sig högst upp på ordförandeskapets dagordning .
Genom att besvara de frågor som Ana Terrón i Cusí har ställt , skall jag försöka besvara de som handlar om inrikes frågor , och min kollega kommer därefter att ta upp de rättsliga frågorna .
Som ni känner till tillämpas Schengenregelverket helt i tio länder , och under år 2000 kommer arbete att bedrivas för att Schengenregelverket skall kunna träda i kraft i Danmark , Finland och Sverige , liksom i Island och Norge .
Rådets generalsekretariat har offentliggjort en dokumentsamling som innehåller hela Schengenregelverket , och väntar på offentliggörande i EGT när alla översättningar finns tillgängliga .
Denna samling finns för närvarande på sex språk och övriga översättningar är på väg att avslutas .
En annan fråga handlar om programmen för invandring och asyl och tillämpningen av dem i länderna i Central- och Östeuropa .
I mars 1998 antog rådet programmet Odysseus , ett program för utbildning , utbyte och samarbete inom asyl- , invandrings och yttre gränskontroll .
Det tillämpas i unionens femton medlemsstater och förutser möjligheten att associera ansökarländerna liksom eventuellt tredje land .
Programmet täcker perioden 1998 till 2002 och det beräknade beloppet för dess genomförande är 12 miljoner euro .
Ansökarländerna kan associeras till projekt som förvaltningskommittén valt ut och som har samband med programmets mål .
Anslagsbeloppet för 2000 är beräknat till tre miljoner euro .
Inom ramen för programmet 1999 fick kommissionen 80 ansökningar om ekonomiska medel till ett totalt belopp på 7,5 miljoner euro , medan det disponibla anslagsbeloppet för 1999 är 3 miljoner euro .
Kommissionen föreslog att behålla 35 projekt , av vilka 12 på 50 000 euro och 23 på mer än 50 000 euro .
När det gäller Oisin-programmet för budgetåret 1997 , antogs projekt som innehöll seminarier , utbildning , utbyte mellan tjänstemän , undersökningar och studier och verksamhet av operativ karaktär .
Av 62 projekt omfattade 7 ansökarländer .
När det gäller Schengeninformationssystemet ( SIS ) kan vi här säga att medlemsstaterna anser den verksamheten och användningen av SIS som mycket positivt .
Det ökade antal positiva resultat visar på effektiviteten i systemet och antalet signaler upphör inte att öka .
För att utveckla tullinformationssystemet uppnåddes ett avtal med kommissionens avdelningar om ett system som gör det möjligt att arbeta med en provisorisk tillämpning av konventionen om tullinformationssystem så snart ett visst antal ratifikationer av denna konvention har gjorts .
Sedan talade ledamoten om ett interinstitutionellt avtal .
Jag borde ta upp denna sista punkt efter min kollega från justitiedepartementet , men det jag kommer att säga kommer givetvis från ett utbyte av intryck i rådet , och framför allt mellan oss två .
Förutom det jag redan har tagit upp tidigare , det vill säga , en ny relation med kommissionen och parlamentet för en tätare förbindelse där parlamentet informeras i tid angående de frågor som rådet kommer att diskutera , skulle jag här inför er vilja uttrycka vår beslutsamhet att rådgöra med Europaparlamentet , inte bara i de fall som fördraget föreskriver , för det är vi tvingade till , utan också att informera och rådgöra med parlamentet när vi anser det viktigt att utvidga denna typ av samråd , och i direkt kontakt med kommissionen , om den anser att parlamentet bör yttra sig i denna fråga .
När det gäller informationen kommer vi att kommunicera med parlamentet om alla de områden som är viktiga för skapandet av ett område med frihet , säkerhet och rättvisa , så att det blir möjligt för detta partnerskap mellan rådet och parlamentet , grundat i kommissionen och på det utmärkta arbetet av kommissionär António Vitorino som alltid är så framåt , att göra det portugisiska ordförandeskapet till en riktpunkt i skapandet av ett område med frihet , säkerhet och rättvisa .
( Ihållande applåder ) Herr talman , mina damer och herrar , herr kommissionär !
Då jag inte har varit ledamot i Europaparlamentet tidigare förstår ni nog att min sinnesrörelse över att vara närvarande här är större än den som min kollega Fernando Gomes känner .
Som ledamoten Anna Terrón sade i sitt inlägg präglas år 1999 av en dominans för de rättsliga och inrikes frågorna , ett år av stora förväntningar .
Förväntningar som konkretiserades genom att Amsterdamfördraget trädde i kraft , förväntningar som konkretiserades i slutsatserna från rådet i Tammerfors , men förväntningar som det är viktigt att i år överföra i konkret handling , att genomföra , och därför är vi alla medvetna om att det är viktigt att rådet så snabbt som möjligt kan godkänna den resultattavla som kommissionär António Vitorino har i uppdrag att genomföra .
Jag måste än en gång uttrycka vår djupa önskan om att det portugisiska ordförandeskapet skall kunna avsluta det politiska avtalet om en resultattavla under det informella rådet i Lissabon den 3 och 4 mars .
När det gäller de konkreta frågor som ledamoten Anna Térron ställde , skulle jag vilja dela in dem i tre grundläggande ämnen : kampen mot den organiserade brottsligheten , det rättsliga nätverkets verksamhet , särskilt i straffrättsliga frågor , och frågor gällande Europol .
När det gäller kampen mot den organiserade brottsligheten , innebar år 1999 förverkligandet av några viktiga åtgärder från handlingsplanen i Wien , främst det som ledde till undertecknandet av stadgan för europeiska yrkesorganisationer och utvecklingen av samarbetet och etablerandet av kontaktpunkter mellan medlemsstaterna angående viktigt informationsutbyte i kampen mot penningtvätt ; jag vill också peka på det finländska ordförandeskapets initiativ vad gäller ett beslut i rådet som nu behandlas i den blandade gruppen .
Detta är ett område där vi måste fortsätta att fördjupa arbetet , inte bara för att få igenom unionens strategi i kampen mot den organiserade brottsligheten under det nya årtusendet , utan också för att ta oss förbi de svårigheter som härrör från det existerande lappverket , framför allt på rådsnivå , i bedömningen av hur kampen mot den organiserade brottsligheten skall ske , och i denna mening , vill jag understryka vikten av att vi bidrar till det samarbete vi håller på att utveckla tillsammans med det franska ordförandeskapet , för att genomföra ett RIF-Ekofin " jumboråd " som , för att det inte bara skall ebba ut i en ren massmediahändelse , bör föregås av ett noggrant förberedelsearbete baserat på en blandad kommitté vars sammansättning det portugisiska ordförandeskapet redan har lagt ett förslag om .
En annan viktig fråga i samband med kampen mot organiserad brottslighet handlar om förbindelserna med tredje land .
Här är det viktigt att det går att utarbeta en gemensam handlingsplan , förutom det arbete som bedrivs i expertgruppen om avtal inför anslutningen , mellan Europeiska unionen och Ryska federationen för att bekämpa den organiserade brottsligheten , vilket befinner sig i en avslutningsfas , liksom att genomföra officiella möten med medlemsstaters tjänstemän i Moskva , och utveckla en samling andra initiativ .
Det finns ett område som handlar om unionens ingripande inom ramen för FN-konventionen och respektive protokoll mot den organiserade brottsligheten och de konventioner som har utformats inom ramen för Europarådet , främst om " cyberbrottsligheten " .
Då det handlar om en fråga som har fått en viktig plats inom programmet för rättsliga och inrikes frågor , anser ordförandeskapet det vara av intresse att , i ljuset av principerna i avdelning VI i fördraget , finna lämpliga former för att förse Europaparlamentet med bättre information om hur dessa förhandlingar går och vad de resulterar i , inom ramen för FN-konventionen .
När det handlar om det rättsliga nätverket , har ett viktigt arbete utförts , främst genom igångsättandet av verksamheten , i slutet av 1999 , för det europeiska rättsliga nätverkets telekommunikationssystem , och inom ramen för den blandade gruppen utvecklades en samling åtgärder för genomförandet av handlingsplanen från 1997 .
Men vi understryker att det är viktigt att så snart som möjligt , godkänna strategin för det nya årtusendet så att det arbete som har bedrivits inom ramen för den tidigare handlingsplanen får ny skjuts och kan fortsätta .
Även beträffande det rättsliga samarbetet , har viktiga steg tagits när det gäller det straffrättsliga skyddet för euron och ett rambeslut befinner sig i Europaparlamentet för rådfrågning , ett rambeslut som är av mycket viktig strategisk betydelse .
Vi anser att det straffrättsliga skyddet av euron kräver att vi undviker en mängd instrument och att vi därför måste anstränga oss gemensamt för att i mars kunna godkänna ett enda instrument som gemensamt behandlar de frågor som skall behandlas , dels de som består av initiativ som redan har lagts fram av Frankrike , dels de som kommissionen själv har betonat att det är viktigt att anta .
Det är viktigt att på detta område genomföra åtgärder när det gäller ett ömsesidigt erkännande av rättsliga beslut och vi anser att det är möjligt genom det arbete som redan har bedrivit att åtminstone beträffande konfiskering av tillgångar , inom kort vidtar åtgärder som gör ett ömsesidigt erkännande av besluten möjligt .
Slutligen , när det gäller Europol , som inledde sin faktiska verksamhet under just 1999 , vilket fick rådet att godkänna en rad instrument , som parlamentet känner till , för att få i gång verksamheten i Europol , kvarstår tydligtvis en grundläggande fråga som handlar om den demokratiska och den rättsliga kontrollen av Europol , frågor som givetvis får en annan dimension genom det politiska ställningstagandet i Tammerfors om att fördjupa Europols befogenheter och framför allt att ge den en operativ dimension .
Det franska ordförandeskapet gav oss ett viktigt arbetsdokument med olika scenarier för att möta och lösa frågorna om demokratisk och rättslig kontroll av Europol .
Det portugisiska ordförandeskapet kommer inom kort att ta initiativ till ett arbetsdokument om nätverket Eurojust , för även om det inte är helt nödvändigt att den rättsliga kontrollen av Europol utövas av Eurojust , kan vi inte nu utesluta att det kan vara ett alternativ .
Det är därför viktigt att den debatt som rådet håller om utvecklingen av Europol och Eurojust sker samtidigt för att vi skall kunna fatta besluten samtidigt .
Jag anser att det är inom denna ram , och inom ramen för den dialog rådet och parlamentet måste skapa om utvecklingen av Europol och Eurojust , som vi får möjlighet att finna en godtagbar institutionell lösning för förbindelserna mellan rådet och parlamentet när det gäller Europol .
Vi känner till parlamentets ståndpunkter och vi vet att parlamentet känner till rådets rättstjänsts ståndpunkter .
Jag tror att det är genom att lösa frågan om den demokratiska kontrollen av Europol som denna fråga kommer att få en definitiv lösning och en lösning som mobiliserar och stärker det institutionella samarbetet mellan alla .
( Applåder ) Herr talman !
Mina damer och herrar , ärade rådsmedlemmar !
För det första , utan att gå in på någon tävling om känslor med ministrarna , vill jag säga att jag inte känner sinnesrörelse , jag känner mig förvirrad av att i ordförandeskapet för första gången ha två personliga vänner och jag hoppas att detta faktum inte kommer att förändra maktdelningen , som är viktig för vår union .
Sedan skulle jag vilja gratulera ledamoten Anna Terrón till att ha tagit upp den fråga som gett upphov till den första debatten i år under denna mandatperiod om skapandet av ett område med frihet , säkerhet och rättvisa , samt tacka alla ledamöter som i de olika utskotten har deltagit aktivt i förberedandet av denna debatt , liksom företrädarna för de nationella parlamenten och det civila samhället .
Jag vill i detta första inlägg ge parlamentet kommissionens syn på det mest betydelsefulla som hände under år 1999 .
Jag tycker att jag med övertygelse , men också med tillfredsställelse , kan säga att år 1999 var en vändpunkt och ett befästande av unionen i frågorna om frihet , säkerhet och rättvisa .
Det har redan sagts här att Amsterdamfördraget trädde i kraft i maj , och detta parlament ansåg att den mest långtgående nyheten i detta fördrag var erkännandet av att det var nödvändigt att skapa ett område med frihet , säkerhet och rättvisa .
Detta utgör samtidigt ett kvalitativt mycket viktigt hopp framåt och ett logiskt och oumbärligt steg i unionens utveckling , efter skapandet av den inre marknaden , införandet av den gemensamma valutan och lanserandet av en gemensam utrikes- och säkerhetspolitik .
Detta projekt är , mer än ett institutionsprojekt , ett projekt för medborgarna i vår gemensamma union .
Därför måste alla medborgare i unionen få en verkligt fri rörlighet , och vi måste erkänna att denna bara är meningsfull om den genomförs i ett säkert sammanhang , med stabil grund i ett effektivt rättsligt system som alla har tillgång till under enkla och lika förutsättningar , och som medborgarna kan lita på .
Unionens ansträngningar att förverkliga ett område med frihet , säkerhet och rättvisa befästes i Tammerfors .
Jag skulle vilja understryka det starka politiska budskap som Europeiska rådet gav , där det framhöll den betydelse stats- och regeringscheferna lade vid ett viktigt förslag , liksom vid antalet politiska riktlinjer och prioriteringar som kommer att göra detta område verkligt , enligt en progressiv strategi , inom ett femårigt perspektiv och detta område har framför allt tre beståndsdelar : Frihet , säkerhet och rättvisa .
År 1999 präglades också av det tyska ordförandeskapets initiativ att utarbeta en stadga om grundläggande rättigheter i unionen .
I Europeiska unionens nuvarande utvecklingsfas , anser jag att det vore lämpligt att samla de gällande grundläggande rättigheterna på unionsnivå i en stadga , för att göra dem mer synliga och tillgängliga för alla medborgare .
Som jag redan har sagt flera gånger så är jag för , och kommissionen är för , att utarbeta en stadga som , grundad på en dynamisk process , återspeglar medlemsstaternas gemensamma konstitutionella traditioner och de allmänna principerna i gemenskapsrätten , och inte bara reducerar dem till en formulering med minsta gemensamma nämnare .
Som företrädare för kommissionen kommer jag att vaka över att stadgan och dess åtgärder befäster en union , som grundas på en rad grundläggande rättigheter som är en del av Europas gemensamma arv .
Bara så kan vi bidra till att legitimera utvidgningsprojektet av unionen i alla europeiska medborgares ögon , en utvidgning som grundas på respekten för rättigheter och friheter , en garanti för människors och egendoms säkerhet och med ett effektivt rättsligt skydd , det vill säga , en union som är grundad på politiska värden som de nuvarande demokratierna bygger på .
Jag tänker inte utelämna att 1999 också var det år då mandatperioden 1999-2004 inleddes i Europaparlamentet och den nya kommissionen tillträde och därmed en kommissionär med exklusivt ansvar för det rättsliga och inrikes området .
Förutom dessa händelser , skulle jag vilja påminna parlamentet om några saker som antogs under år 1999 .
Kommissionen lade fram ett förslag till förordning i fråga om invandring , gränser och asyl , för skapandet av databasen " Eurodac " , förslaget till direktiv om villkoren för tredjelandsmedborgares inresa och vistelse i unionens medlemsstater för att återsamla familjer , inom ramen för en bestämd integrationspolitik av dem som vistas legalt i unionen .
Vi satte i gång en debatt om ett meddelande om gemensamma förfaranden angående asyl och en rekommendation till beslut som bemyndigar kommissionen att förhandla om ett avtal med Island och Norge om en utsträckning av de bestämmelser som Europeiska unionens medlemsstater tillämpar enligt Dublinkonventionen till dessa båda länder .
Kommissionen bidrog aktivt till arbetet i högnivågruppen om asyl och invandring och slutligen , i december , lade den fram ett förslag till skapandet av europeiska flyktingfonden .
På området för rättsligt samarbete lade kommissionen fram förslag till förordningar för att göra vissa konventioner till gemenskapsfrågor : om rättsligt samarbete och verkställighet av domar av civil eller kommersiell natur , ( Bryssel-I ) ; en annan , angående erkännande och verkställighet av domar i äktenskapsmål ( Bryssel-II ) och ännu en annan , delgivning i medlemsstaterna av handlingar i mål och ärenden av civil eller kommersiell natur .
Vi lade också 1999 fram ett meddelande om brottsoffer i unionen och inledde därigenom en diskussion som i Tammerfors tog ett steg framåt och som innehåller krav på minimibestämmelser om skydd för brottsoffer , speciellt tillgång till rättslig hjälp och rätt till ersättning för skador , inklusive rättsliga kostnader .
Jag vill också nämna förslaget till beslut om åtgärder för att bekämpa bedrägeri och förfalskning som rör andra betalningsmedel än kontanter .
Inom ramen för unionens lagstiftning om ekonomisk brottslighet , lade kommissionen fram ett förslag till revidering av direktivet om penningtvätt .
Vi deltog 1999 i starten av Europol , och från kommissionen hoppas vi uppriktigt , särskilt efter vad det portugisiska ordförandeskapet sade här i dag , att den nya perioden för rättsliga och inrikes frågor , och de påbörjade diskussionerna om att införa nya befogenheter för Europol i Amsterdamfördraget , också skall följas av en diskussion om demokratisk kontroll och förbindelserna mellan Europol och behöriga rättslig instans , nämligen Eurojust .
Kommissionen lade 1999 även fram sitt bidrag till en europeisk handlingsplan för narkotikabekämpning , vilken ligger till grund för den strategi som godkändes av Europeiska rådet i Helsingfors .
Denna åtgärdslista , som inte är uttömd , har bidragit till att jag i dag , inför rådets ordförandeskap och ledamöterna , med stor övertygelse kan säga att , om 1999 var ett år som befäste unionens verksamhet inom detta grundläggande område så hoppas jag också att 1999 innebär början på en ny period , en strävan att skynda på skapandet av ett område med frihet , säkerhet och rättvisa .
Därför kommer år 2000 utan tvivel att bli ett år för att pröva hur de europeiska institutionerna klarar att möta medborgarnas krav om fri rörlighet , i respekten för rättigheter och i garantier för säkerhet och stabilitet , genom ett adekvat rättsligt skydd .
Vi kan också säga att år 2000 för rådet , parlamentet och kommissionen kommer att vara ett prövoår för den politiska viljan att ta Amsterdam på allvar och lägga grunden för en utvidgad politisk union under nästa decennium .
Som jag har sagt är kommissionen medveten om sin del av ansvaret och i detta sammanhang har den snart avslutat ett första utkast till förslag till resultatöversikt , en scoreboard , där alla institutioner och andra berörda delar kan börja utvärdera de framsteg som skett genom införandet av nödvändiga åtgärder och uppfyllandet av de tidsfrister som fastställts i Amsterdamfördraget , handlingsplanen från Wien och slutsatserna från Tammerfors .
Denna resultatöversikt kommer inte bara att vara ett instrument för programplanering av lagstiftning utan också , och framför allt , ett instrument för att stärka alla europeiska institutioners öppenhet och ansvar inför medborgarna .
Detta därför att det är för medborgarna som vi utvecklar ett område med frihet , säkerhet och rättvisa .
Framstegen beror inte på kommissionen , inte på rådet , inte ens på Europaparlamentet , utan på de europeiska institutionerna i helhet och på medlemsstaterna själva , då vissa uppgifter på resultatöversikten , vilket redan har sagts här , anförtros medlemsstaterna enligt subsidiaritetsprincipen .
De närmaste veckorna kommer jag att genomföra en rundresa i huvudstäderna för att lyssna på ministrarna för rättsliga och inrikes frågor .
Jag räknar med att debattera projektet med resultatöversikt med Europaparlamentet och med det civila samhället .
Vi räknar med att efter dessa konsultationer lägga fram slutversionen inför rådet för justitie- och inrikesministrar , under det portugisiska ordförandeskapet .
Min avsikt är att denna resultatöversikt skall bli ett instrument för politisk och strategisk inriktning för alla institutioner men också ett instrument för opinionsundersökningar .
Därför inser jag - och det är en utmaning som jag tror att vi alla ställs inför - , att utveckla en kommunikationsstrategi som kan göra det mervärde som unionen innebär för allmänheten i dess dagliga liv , tillgängligt och begripligt i dessa viktiga områden för medborgarna , i respekten för lagligheten och i grunden själva demokratin .
Förutom resultatöversikten skulle jag vilja nämna att kommissionen räknar med att under år 2000 lägga fram följande initiativ - och jag skulle här vilja understryka att jag gratulerar till att det portugisiska ordförandeskapet betraktar utvecklingen av detta område som en av sina prioriteringar i arbetsprogrammet .
Jag hoppas att det blir möjligt , under det portugisiska ordförandeskapet , att tydligt utveckla en interinstitutionell samarbetsanda , vilket också är det politiska budskapet från Tammerfors , och att denna interinstitutionella samarbetsanda följs upp av de efterföljande ordförandeskapen .
När det gäller invandring och asyl , räknar kommissionen med att kunna lägga fram förslag till utformningen av ett gemenskapsinstrument för tillfälligt skydd av flyktingar ; inleda analysen av kriterier och villkor för att förbättra genomförandet av Dublinkonventionen och ett övervägande att förändra dess rättsliga grund i enlighet med Amsterdamfördraget ; fortsätta debatten utifrån det meddelande som redan har spridits om bestämmelser som leder till ett gemensamt asylförfarande i hela unionen ; och lägga fram lagstiftningsförslag om att bevilja uppehållstillstånd till de offer för människohandel som samarbetar med rättsväsendet mot nätverken för människohandel .
Jag räknar också med att kunna bidra till ett klargörande av handlingsplanernas roll inom arbetet i högnivågruppen om asyl och invandring och gå vidare med antagandet av gemenskapsavtal för återinresa , genom att införa klausuler för detta ändamål .
I en central fråga angående den fria rörligheten såsom resa över de yttre gränserna i medlemsstaterna kommer jag under de närmaste dagarna att lägga fram ett förslag till förordning som förnyar listan över tredje land vars nationaliteter måste ha visering för att kunna passera de yttre gränserna .
Inom det rättsliga samarbetet hoppas jag innerligt att det , förutom ett initiativ om lagen som är tillämplig på förpliktelser ej angivna i kontrakt blir möjligt att lägga fram ett förslag till minimibestämmelser som garanterar en lämplig nivå av rättshjälp över hela unionen vid gränsprocesserna .
Jag räknar också med att kunna fortsätta arbeta med nya gemensamma processregler specifikt för att förenkla och påskynda av gränsöverskridande rättsliga processer i mindre fall gällande handel och konsumenter , matpensioner och ej besvarade åtal .
I uppföljningen av slutsatserna från Tammerfors och Helsingfors kommer kommissionen att lägga fram sitt bidrag till definitionen av en unionens strategi för att förebygga och bekämpa den organiserade brottsligheten .
Vi kommer att organisera och stödja åtgärder och särskilt debatten om behovet att utarbeta ett lagstiftningsprogram för genomförande av principen om ömsesidigt erkännande av domar i straffrätten .
Kommissionen räknar också med att lägga fram specifika åtgärder för förebyggande av brottslighet för att utveckla utbytet av den bästa praxisen på området , speciellt förebyggande av brottslighet i städerna och ungdomsbrottslighet , och lägga fram en rättslig grund för ett program , finansierat av gemenskapen .
Kommissionen kommer också att bidra till ordförandeskapets arbete för att klargöra den rättsliga ramen och den administrativa polisiära och rättsliga samarbetsramen för att bekämpa penningtvätt , i ett perspektiv som i hög grad överskrider gränserna mellan pelarna .
Kommissionen kommer att uppfylla det ansvar den fick i Tammerfors för att lägga fram förslag till antagande av gemensamma definitioner , åtal och sanktioner mot människohandel och ekonomiskt utnyttjande av invandrare och sexuellt utnyttjande av kvinnor och barn , med särskild tonvikt lagd på kampen mot användande av de nya kommunikationsmedlen , främst Internet , för spridning av barnpornografi .
Vi förbereder också ett meddelande för att diskutera medlen för att skapa ett samhälle med säkrare information och kunskap och för att kunna bekämpa datorbrottslighet .
År 2000 innebär också inledningen av tillämpningen av den europeiska strategin mot narkotika för perioden 2000-2004 .
Kommissionen kommer på detta område och i samarbete med det portugisiska ordförandeskapet och Europaparlamentet , att ge allt sitt stöd till den interinstitutionella konferensen i februari om narkotikaproblematiken .
Beträffande Schengen skulle jag , utan att nu gå in på rådets behörighetsområde , och särskilt när det gäller integreringen av Schengenregelverket inom gemenskapsramen , vilja understryka att kommissionen , i den aktuella frågan om återupprättandet av gränskontroll , än en gång upprepar sin beredskap att fördjupa formerna för en bättre kontroll av tillämpningen av artikel 2.2 i Schengenkonventionen , så att den blir mer tvingande .
Återinrättandet av viss intern gränskontroll nyligen får mig att dra slutsatsen att det är nödvändigt att göra en detaljanalys av förutsättningarna för att anta ett lagstiftningsinstrument grundat på artikel 62 i fördraget .
Så som betonades i Tammerfors , och med tanke på förberedelserna av Europeiska rådet i Feira , i juni 2000 , måste vi sammanfatta innebörden av den nya externa dimensionen i de inrikes och rättsliga frågorna med perspektiv på ett antagande av politiska strategier mellan pelarna för att förstärka sammanhållningen i unionens inrikes- och utrikespolitiska förbindelser för att bidra till att befästa unionen i världen .
Jag vill emellertid understryka att alla dessa åtgärder givetvis måste ske med hänsyn till de principer som beslutats vid Europeiska rådet i Helsingfors i förhållande till ansökarländerna , så att dessa ansökarländer samarbetar och så snart som möjligt knyts till projektet att skapa ett område med frihet , säkerhet och rättvisa .
Det är för övrigt viktigt att komma ihåg att förhandlingarna om rättsliga och inrikes frågor inleds år 2000 med den första gruppen ansökarländer och jag hoppas att vi skall kunna göra stora framsteg i förberedelserna av de förhandlingsärenden angående den andra gruppen som i Helsingfors godkändes för anslutning .
Slutligen skulle jag vilja säga att kommissionen försöker vara i en pole position i presentationen av förslag för att kunna följa upp genomförandet av Amsterdamfördraget .
Jag hoppas att kommissionen och rådet kommer fram till ett avtal om delat ansvar i utövandet av initiativrätten och ledningen av själva lagstiftningsprocessen .
Som jag sade till parlamentet , den uppgift vi har framför oss är enorm och ambitiös , kommissionen behöver vara utrustad med nödvändiga mänskliga resurser för att kunna möta denna utmaning och hoppas få parlamentets stöd , och varför inte rådets , för att garantera dessa resurser och mål , så att skapandet av ett område med frihet , säkerhet och rättvisa i unionen blir verklighet så snart som möjligt och på så sätt kan vi alla bidra , i en anda av interinstitutionellt samarbete , för att genomföra detta projekt , vilket utan tvivel är " kronjuvelen " i Amsterdamfördraget .
Herr talman , ärade kolleger !
Efter att denna församling under 40 år ägnat sig huvudsakligen åt att etablera en gemensam inre marknad har vi nu en ny stor uppgift i att skapa ett område av frihet , säkerhet och rätt .
Det är en uppgift som vi emellertid endast kommer att kunna lösa framgångsrikt om alla unionens institutioner arbetar gemensamt med ömsesidig respekt mot det ambitiösa målet , under beaktande av respektive befogenhetsområden .
Kommissionär Vitorino , medan jag vill beteckna samarbetet med er som harmoniskt och fruktbart så har jag ofta saknat ord för att beskriva det uppträdande som rådet visat prov på i förbindelserna med oss .
Det har verkat - som kollegan Schulz en gång träffande sagt i utskottet - som om rådet under området av frihet , säkerhet och rätt tänkt sig ett område för egen oansvarighet , för säkerhet att inför parlamentet och rätten göra och låta ske enligt eget godtycke .
Herr minister Gomes , jag har förstås uppfattat era redogörelser om detta .
Följaktligen hoppas jag på en tydlig förbättring i samarbetet under det portugisiska rådsordförandeskapet .
Jag vill lyfta fram tre punkter vilka för oss medlemmar i Europeiska folkpartiets grupp måste vara tyngdpunkter i skapandet av ett sådant område .
För det första : uppbyggandet av en gemensam asylrätt och en fördelning av de bördor som uppkommer i samband med mottagande av flyktingar .
Först måste rådet äntligen tillse att Eurodac blir utfärdat för att skapa en grundförutsättning för fördelning av asylsökandena .
Vad beträffar en asylrätt som gäller över hela Europa har förvisso ett par ansatser blivit synliga genom Wien och Tammerfors .
Dessa ansatser visar emellertid dessvärre snarare på de svårigheter som finns i stället för att komma med lösningsförslag .
Företrädarna i rådet uppmanas därför att blicka ut över sina egna nationella murar och skapa ett enhetligt asylförfarande för hela unionen .
Det kan heller inte vara riktigt att några få hjälpvilliga medlemsländer skall tvingas bära hela bördan av flyktingeländet på vår kontinent .
En överenskommelse om en fördelning av bördorna måste av den anledningen ha högsta prioritet .
För det andra : utbyggnaden av ett alleuropeiskt bekämpande av den organiserade brottsligheten , bland annat via Europol och Eurojust .
Det planerade inrättandet av Eurojust framstår för oss som ett viktigt framsteg från Tammerfors som nu måste genomföras snarast .
Vi välkomnar det faktum att Europol till slut har kunnat påbörja sitt arbete .
Rådet får dock ej bortse från att det för att effektivisera brottsbekämpningen inte räcker med den i Tammerfors beslutade fördelningen av Europols uppgifter , utan att det måste ingå såväl en personell förstärkning som en uppgiftsfördelning ända ned till den operativa nivån .
Det är inte så att vi ropar efter ökad kontroll och mer kontroll över själva Europol ; för oss gäller här snarare talesättet : " Mindre är ibland mer ! "
Om en huvuddel av Europols medarbetare för närvarande framför allt är sysselsatta med att kontrollera sig själva i datasäkerhetsrättsligt hänseende varvid man inhämtar undersökningar från 15 olika nationella parlament är detta mycket kontroll , men en ineffektiv kontroll .
Vi vill ha mindre virrvarr i kontrollen men ökad parlamentarisk kontroll genom Europaparlamentet , och detta utan att Europols arbete skall hindras .
Samtidigt stöder vi inrättandet av en europeisk polisakademi , vilket föreslagits i Tammerfors , såsom ett steg i rätt riktning .
För det tredje : utvidgningen av parlamentets rättigheter i detta sammanhang .
Om det bara blir diplomater och byråkrater som bestämmer över inrättandet av en anordning som medger unionen att även ingripa i de grundläggande fri- och rättigheterna för unionens medborgare , medan de valda företrädarna i Europa inte kan annat än bara följa utvecklingen som kaniner gör med ormens rörelser , så kommer denna anordning aldrig att accepteras av medborgarna .
Det är därför på tiden att parlamentet härvidlag tillerkänns medbeslutanderätt och - som redan sagts - att principen om demokratisk kontroll stärks .
Vi vill ha ett område av frihet , säkerhet och rätt för medborgarna i Europa och inte mot dem .
Högt ärade herr talman , mina kära kolleger !
Jag behöver inte säga något mer om rådet .
Föregående talare har redan gjort det med hjälp av ett citat av mig från det senaste utskottssammanträdet .
Varför har rådet ett sådant motstånd mot att samarbeta med oss i uppbyggnaden av området av säkerhet , frihet och rättvisa ?
Den frågan kommer ständigt för mig .
Jag vill försöka belysa den en smula som jag ser Byggandet av ett område för säkerhet , frihet och rättvisa beror skiljelinjen mellan den nationella suveränitetens grundläggande delar .
Polis och rättsväsende är två väldefinierade delar som ingår i självstyret ; dvs. detta är känsliga politikområden i medlemsländerna - det börjar närma sig ett överförande av politikområden till gemenskapen , alltså ett delegerande av befogenhet från den nationella huvudstaden , t.ex.
Lissabon , Berlin eller Paris till Bryssel .
Det är ett stycke överföring av makt .
Det är självklart att det är mycket , mycket svårt att skiljas från förmedlade , traderade verkställighetsformer också när man själv inser att ett polisiärt samarbete är nödvändigt ; den internationella brottsligheten kan bara bekämpas på Europanivå .
Då är det nödvändigt att dra konsekvensen av det och säga : Vi måste då också överföra instrumenten organisatoriskt och juridiskt till gemenskapen .
Det innebär att de regeringar som skall göra det och inser nödvändigheten av det på samma gång inser att de i och med förverkligandet också beskär sin egen makt .
Dessutom finns det ett Europaparlamentet med mycket komplex funktion .
Men någon gång måste vi hitta en lösning på problemet .
Ty om vi fortsätter på samma sätt som vi gjort hittills kommer följande att inträffa : Säkerhetsdebatten , debatten om medborgarnas rättigheter marginaliseras i de nationella parlamenten genom konstruktionen av till hälften nationell och till hälften europeisk uppbyggnad .
Debatten når inte ända fram till Europaparlamentet , medan rådet sammanträder bakom lyckta dörrar .
Om uppbyggnaden av området av säkerhet , frihet och rätt förblir en hemlig anordning kan vi inte vinna medborgarnas gillande av den bakomliggande idén .
Dvs. när vi diskuterar detta handlar det om demokratins stabilitet .
Det är därför som jag blir så upprörd - alltså inte över ministerrådet .
Ministrarna är i regel valda ledamöter .
Kollegan Gomes , kollegan Costa , kollegan Vitorino , vi har allihopa i princip samma bakgrund .
Jag vill emellertid rikta en vädjan till rådets byråkrati .
Följande princip gäller : Den som förbereder beslut - och det gör rådets byråkrati , den föregriper dem - bör nog visa litet mer demokratiskt mod .
( Applåder ) Jag vill bara helt kort nämna ytterligare en aspekt , jag har ju inte mycket tid kvar .
Scoreboard , på tyska låter det som skateboard .
Jag säger därför att vi behöver en tidsplan som anger vilka frågor som skall förverkligas när och av vem .
Vitorino-planen - att genomföra tydligt preciserade projekt på en tydligt definierad tid - är vad vi behöver .
Detta förmår kollegan Vitorino , som jag vill tacka för hans anförande , enbart under förutsättning att han får de nödvändiga finansiella och personella resurserna .
Låt oss ge honom dem , så att han kan göra snabba framsteg vilket gynnar oss alla .
Jag välkomnar varmt det faktum att det portugisiska ordförandeskapet sätter rättsliga och inrikes frågor högt , om inte högst , på prioriteringslistan .
Jag blev också glad att höra kommissionär Pattens kommentarer i förmiddags om en fond för snabba åtgärder vid säkerhetskriser .
Kanske detta kan få slut på skandaler som misslyckandet med att sätta in den utlovade polisstyrkan i Kosovo .
Låt mig bara betona tre områden bland många där vi behöver se snabba framsteg .
Det första rör asyl .
Det är nödvändigt att upprätta ett gemensamt europeiskt system , men det skall grundas på rättvisa , fullständig respekt för Genèvekonventionen och anständiga mottagningsförhållanden , inklusive ett slut på de rutinmässiga kvarhållandena .
Ett asylbeslut bör kunna fattas inom några månader - inte inom några år .
Det andra området rör frihet : Frihet att flytta och bosätta sig var man vill inom unionen ; informationsfrihet ; frihet att rösta på alla som har ett europeiskt medborgarskap - och detta omfattar inte bara medborgare i medlemsstaterna , utan även medborgare från tredje land .
Låt våra medborgare få veta att vår gemensamma politik rörande rättsliga och inrikes frågor handlar om frihet , inte bara om förtryck .
Det sista området jag vill nämna handlar om konvergering av civil- och straffrättsliga system .
Euroskeptikerna hävdar att detta är ett hot mot suveräniteten , slutet för nationalstaten , osv. men fallet som rör den misstänkte som var efterlyst för utfrågning i samband med morden på tre kvinnor i Frankrike , inklusive den brittiska studentskan Isabel Peake , som blev avslängd från ett tåg , visar varför vi behöver ett ömsesidigt erkännande .
Mannen som arresterades och släpptes i Madrid , har nu blivit utlämnad efter att ha suttit arresterad i Lissabon .
Vad euroskeptikerna än säger ligger det i allas vårt intresse att det sker ett samarbete kring sådana frågor .
Sammanfattningsvis , som redan nämnts , är det nödvändigt - och jag hoppas att detta tas upp på regeringskonferensen - att det ändras till medbeslutandeförfarandet inom dessa områden , med demokratisk och rättslig granskning .
Herr talman , angående år 1999 kan jag bara säga följande helt kort : Efter den finska kylan är Portugals solsken hjärtligt välkommet .
Jag hoppas att det också går bra .
En för Europa viktig händelse under 1999 när det gäller området av frihet , säkerhet och rättvisa var helt säkert toppmötet i Tammerfors .
Men fortfarande kvarstår åtskilliga frågor att besvara .
Många svar väntar vi ännu på .
Dock efter Tammerfors har vi fått en obalans mellan de positiva åtgärder som faktiskt vidtogs och rena avsiktsförklaringar .
Det återstår fortfarande att besluta om medborgarskapsregleringen samt om integrationen av människor från tredje land .
Å andra sidan har man nu tagit initiativ till högst konkreta åtgärder på temat säkerhet .
Framtagandet av en stadga med grundläggande fri- och rättigheter torde bli ett av de stora projekten i den nära framtiden .
När jag tänker på de människor som för närvarande ej är unionsmedborgare känns det dock svårt att förutsäga hur denna stadga kommer att se ut rent innehållsmässigt och vilken utformning i rättslig mening förverkligandet av den kommer att få .
Europolavtalet har nu officiellt trätt i kraft .
Vid mötet i Tammerfors siktade man på att också fördela de operativa befogenheterna .
Men vi kräver alltjämt en revidering av avtalet , vilket syftar till att åstadkomma förbättrade parlamentariska och rättsliga kontrollmöjligheter .
Också vad gäller Eurodac bör avtalet ställas under kritisk belysning .
Parlamentet har modifierat fördragstexten .
Det måste garanteras att rådet går på samma linje som parlamentet .
Vad gäller övriga ämnen har det tyvärr ännu inte tagits några initiativ .
Vi väntar för ögonblicket på det .
Europa såsom ett område av frihet , säkerhet och rättvisa är fortfarande en anordning utan klar reglering på centrala områden .
Vi är dock skyldiga de europeiska medborgarna detta .
Efter att ha hört inrikesministern och justitieministern tala är jag numera optimistisk .
Jag utgår ifrån att vi kommer att lyckas med detta under de kommande sex månaderna .
Herr talman , herr kommissionär , kära kolleger !
Jag tror att den muntliga frågan från Terrón i Cusí är intressant så till vida att den är ett tramp i klaveret , för sex månader efter att vårt nya parlament inrättats måste vi kunna ge ett starkt politiskt budskap till Europas medborgare .
Jag tror att det portugisiska ordförandeskapet positivt kan bidra till det .
Vi känner i dag alla till de ofantliga förväntningarna från våra landsmän när det gäller frihet , säkerhet och rättvisa , bl.a. på det sociala området .
Men deras brist på intresse , deras distans och ibland t.o.m. avsky för politiken tvingar oss att vidta konkreta åtgärder mot svårigheterna .
Det är ett oeftergivligt villkor för att de på nytt skall komma överens med politiken .
För att Europa skall bli en symbol för fred och broderskap måste vi bedriva en djärv och generös politik och hjälpa de sämst lottade .
En verklig handlingsplan mot arbetslösheten måste inrättas , för det är utifrån denna farsot som rasism , främlingsfientlighet , nationalism och den rasistiska extremhögern frodas .
Bland de sämst lottade , och det är viktigt att jag nämner den punkten , har vi invandrarna och flyktingarna .
Villkoren för att praktiskt taget systematiskt kvarhålla och kriminalisera asylsökande är inte längre godtagbara .
Alla asylsökande måste få rätt att höras rättvist och ha rätt till suspensiv talan .
Jag blev av en tillfällighet vittne till en scen med sällsynt våld i förra veckan på Roissys flygplats , där två unga kvinnor , säkerligen illegala invandrare , återfördes till Conakry .
De behandlades som de värsta brottslingar .
De var nakna , släpades i håret över golvet och omringades av en hord kravallpoliser .
Det portugisiska ordförandeskapet måste få ett stopp på detta slag av barbariska vanor .
Vår roll är i stället att åtfölja , garantera , hjälpa dem som flyr från diktaturer .
Kommissionen föreslog att en europeisk fond för flyktingar skulle inrättas .
Parlamentet är mycket positivt till det .
I stället för att komma med undanflykter när det gäller den budget som beviljats fonden tror jag ni kan fatta beslutet att inrätta den .
Ordförandeskapet och rådet kan konkretisera det som förkastats som obegripligt i Tammerfors , även om Tammerfors utgjorde en viktig grund .
På samma sätt kan vi inte nöja oss med att konstatera att de främlingsfientliga strömningarna ökar i Europa och att man banaliserar diskriminering , utan att vidta omfattande åtgärder .
Det krävs harmonisering av lagstiftningen mot rasism .
Vilken inriktning vill ni ge artikel 13 i fördraget ?
Vad tänker ni göra för att främja lika lön för män och kvinnor ?
Hur tänker ni arbeta för att utrota homofobin , rasismen och sexismen ?
Vi måste använda de bästa tillämpningarna från varje land i unionen .
När sex europeiska länder beviljar rösträtt kan er president tillåta sig att utvidga denna rösträtt och valbarhet i de kommunala och europeiska valen till samtliga medborgare från länder utanför unionen , som sedan fem år bor på europeiskt territorium .
Att ge de personer som inte har några identitetshandlingar uppehållstillstånd i vissa länder , däribland ert , måste bli ett exempel för de övriga , för denna grupp utan identitetshandlingar består i dag av sköra människor som befinner sig i händerna på utsugare och som utnyttjas som arbetskraft , vilket gör dem till den moderna tidens slavar .
Rent allmänt måste detta ordförandeskap inleda förändringar när det gäller uppträdande och förhållanden bland våra landsmän tillsammans med minoriteter och invandrare .
Immigrationen är alltför ofta synonym med osäkerhet och våld och rent repressiva lösningar .
Hur skall ni få våra landsmän att förstå att immigrationen i dag , liksom alltid , är en källa till social och kulturell rikedom , vars roll är och förblir nödvändig i vår demografiska miljö .
Vilka åtgärder avser ni att vidta för att uppvärdera invandrarnas plats i samhället och garantera ett verkligt skydd för asylsökande ?
Herr talman !
Det råder stor brist på öppenhet inom området säkerhet , frihet och rättvisa .
Europeiska unionen är en ekonomisk jätte , men vi har inte rätt att spela ofelbara när det gäller vår behandling av flyktingar .
Nivån på rasismen i vårt samhälle är skrämmande .
Under flera generationer skickade Irland iväg sina söner och döttrar till säkra platser över hela världen , men nu när den keltiska tigern skapar ett välstånd som är större än vad vi förväntat oss , visar vi ett mycket fult drag i vår karaktär .
Rasismen i Irland är endemisk .
Det var en ganska stor chock för våra politiska ledare när de förstod att vi nu måste ta en del av de flyktingar som under en lång tidsperiod rest till Europeiska unionen .
Vi har kommit efter när det gäller att ta itu med denna fråga och regeringen gör sitt yttersta för att hinna ikapp .
Viljan finns , men rädslan dröjer sig kvar ; och för att dämpa denna rädsla måste vi hitta ett politiskt och religiöst ledarskap , inte bara i Irland utan över hela Europeiska unionen .
Herr talman !
Vi kan notera att det urskuldande och försiktiga ordförandeskap som under de senaste månaderna har förhindrat en debatt som den vi faktiskt har lyckats genomföra i dag , har upphört .
Jag instämmer till fullo i det som mina kolleger von Boetticher och Schulz sade och anser det vara helt rätt att Europaparlamentet och domstolen måste engagera sig mer i området frihet , säkerhet och rättvisa utan att behöva avstå från sina egna befogenheter .
Men just för att vi inte skall behöva upprepa det spektakel som var sjätte månad urskillningslöst drabbar rådets ordförande , borde kanske detta parlament ha modet att ta ett kraftfullt politiskt initiativ så att nästa regeringskonferens beslutar att genast utvidga medbeslutandet i stället för att vänta i ytterligare fem år .
De två likalydande frågorna som behandlas , bärs fram av ett mantra som numera mer och mer förvandlar politik till en slags ideologi - välklingande , men fördärvlig .
Och våra dagars EU-mantra heter OFSR - område för frihet , säkerhet och rättvisa .
Bakom detta ligger en annan ambition hos kommissionen , rådet och det överväldigande flertalet i denna församling , dvs. att införa ett sådant område .
Och vem stöder då inte säkerhet , frihet och rättvisa ?
Problemet är bara att det inte är något som EU kan införa genom lagstiftning och andra övernationella åtgärder .
Frihet , säkerhet och rättvisa är ett samhälles rotsystem .
Det är en återspegling av varje samhälles historia , dess sociala erfarenheter och politiska utveckling .
Det är inte något som EU kan införa utan att samhället lider skada .
Men det är just här vi hittar det faktiskt rationella i mantrat om säkerhet , frihet och rättvisa .
Uppgiften är inte att säkerställa rättvisa för medborgarna .
Det sker redan genom de nationella rättssystemen .
Uppgiften är att överföra viktiga delar av samhällets straffrätt , kriminalpolitik och rättskipning till EU : s institutioner .
Det handlar om en förstärkt integration som t.o.m. i en bedräglig förpackning innehåller förstärkt repression och kontroll .
Tänk bara på alla åtgärder kring Fästning Europa , Schengen , Eurodac osv .
Varje demokrat hittar två nyckelproblem .
För det första är de planerade åtgärderna helt orealistiska .
Hur föreställer man sig att EU : s institutioner , som redan lider under en tung arbetsbörda , skall kunna genomföra dessa ambitiösa projekt ?
Tänk på de senaste årens mördande kritik av kommissionens brist på anständighet , etik och ansvar .
Det kommer ju också till direkt uttryck i frågan .
För det andra är projekten belastande - ja , lemlästande - för de nationella demokratierna .
Så länge som EU sysslade med den inre marknaden angrep man bara kroppen .
Nu angriper man själen .
Herr talman !
I dag har det nordirländska folket fått bevittna en underlig , ironisk händelse .
Kommissionär Patten har talat i kammaren och försvarat frihet , säkerhet och rättvisa , och trots detta resulterar den rapport han lagt fram för det brittiska underhuset - vilken har accepterats - i att the Royal Ulster Constabulary och dess reserver försvinner och att nordirländare , både protestanter och katoliker , hamnar i händerna på terrorister .
Terroristerna från IRA har inte lämnat inte några vapen , vilket inte heller de protestantiska terroristerna har gjort , ändå tvingas polisen in i ett läge där de inte har befogenheter att bekämpa terroristerna .
Låt mig ta en titt på siffrorna från den dag avtalet undertecknades .
Under 1998 hade vi 55 mord .
Under 1999 hade vi sju mord och då räknas inte offren för bomben i Omagh med , där 29 dödades och 300 skadades .
Mellan 1998 och 1999 överföll och sköt lojalisterna 123 personer , medan republikanerna överföll och sköt 93 personer .
Antalet åtal som väcktes mot lojalisterna under 1999 uppgick till 193 och motsvarande siffra för republikanerna var 97 .
Sedan januari 2000 har det skett sex överfall med skjutvapen som utförts av lojalisterna och två av republikanerna ; lojalisterna har varit inblandade i sex allvarliga överfall , varav ett resulterade i ytterligare ett mord , samtidigt som republikanerna varit inblandade i fem allvarliga överfall .
Herr talman !
Man måste komma till rätta med situationen - detta kan inte fortsätta .
Herr talman !
Amsterdamfördraget har visat sig vara ett viktigt mål för unionen , och en uppgift som alla parlamentsledamöter , rådet och kommissionen bör åta sig under den här mandatperioden är , såsom nämnts , att skapa området frihet , säkerhet och rättvisa .
Rådet i Tammerfors , motor och upphovsman till denna målsättning , föreslog vissa mål , men fem år för att utveckla avdelning IV i fördraget är för lång tid att vänta för att lösa vissa problem som brådskar .
Min första tanke är att parlamentet inte bör utelämnas från de viktiga beslut som skall fattas i den här frågan och att vår delaktighet i beslutsförfarandet måste garanteras , särskilt när det gäller ett projekt för medborgarna , som kommissionären uttryckte sig så väl .
Min andra tanke är att vi skyndsamt måste anta ett gemensamt system för asyl genom att godkänna gemensamma förfaranden , men framför allt genom att sätta stopp för den förvirring som nu råder mellan emigration av politiska skäl och den berättigade av ekonomiska skäl .
De sist antagna utlänningslagarna i mitt land , Spanien , eller i Belgien , är en larmsignal för att immigrationspolitiken skyndsamt måste införlivas .
Min tredje och sista tanke rör unionens externa åtgärder när det gäller immigration och asyl .
Vi varken får eller kan ge ett intryck av att unionen bara försöker skydda sig från vågen av flyktingar och ekonomiska immigranter .
Vi bör välja samarbetspolitik för utveckling med våra grannar i öst och i Medelhavsområdet , men detta skall göras rigoröst med ekonomiska medel och ett nära samarbete med de offentliga institutioner som samarbetar för att skydda de medborgare som får sina mest grundläggande rättigheter kränkta eller som vill emigrera för att täcka sina grundläggande behov .
Avslutningsvis , när det gäller dokumentet om de grundläggande rättigheterna , så måste Europas medborgare få visualisera sitt medborgarskap .
Det räcker inte med euron eller sysselsättning , inte ens med säkerhet .
De behöver den " europeiska själen " , som en framstående spansk professor en gång sade .
Herr talman !
Till skillnad från vissa andra tidigare talare , vill jag ta upp uttalandena från våra portugisiska ministrar och Vitorino .
Orden som denna trio uttalade lät som musik i våra öron , som Ceyhun sade .
Som med all musik måste det vara en fin sång som är lämpligt instrumenterad .
Många av oss i kammaren ser mycket optimistiskt på de kommande sex månaderna .
Sången som skall spelas kommer att vara en som Europas medborgare skall lyssna på , och de vill höra den rätta sången .
Som beskrivits i eftermiddag kommer det ta lång tid att överrösta vissa av de obehagliga sånger som vi hört under valet till Europaparlamentet och under de senaste månaderna .
Amsterdamfördraget och toppmötet i Tammerfors byggde på detta projekt för ett område med frihet , säkerhet och rättvisa i Europeiska unionen .
Ett område är emellertid oerhört viktigt och denna kammare måste delta i detta , dvs. granskning .
Det finns så mycket lagstiftning - och jag välkomnar verkligen det portugisiska programmet som presenterades för oss i förra veckan - men vi måste vara helt säkra på att det granskats , att personerna i detta parlament och ledamöterna vid de nationella parlamenten och de europeiska medborgarna känner till allt i samband med programmet .
Och vi måste se till att innehållet är genomförbart , lämpligt och relevant för de olika länderna .
Låt mig rikta uppmärksamheten mot vissa aspekter av de resolutioner som vi skall behandla under denna eftermiddag , av vilka det hänvisats till en eller två tidigare .
Jag välkomnar styrningen mot erkännandet av rättsliga system i de olika länderna och samarbetet kring brottslighet .
Detta är ett område som de europeiska medborgarna med glädje kommer att acceptera .
Men kommissionen och rådet måste få veta att det finns många i denna kammare som hyser betänkligheter om t.ex.
Eurodac-systemet .
Vi accepterar rådets dominerande roll i detta sammanhang , men det finns reservationer och jag är säker på att rådet kommer att lyssna på argumentationen från de valda parlamentarikerna när de går igenom saken mer ingående .
Schulz sade tidigare i dag att han inte var säker på vad en " resultattavla " var för något .
Alla som är engelsmän eller britter eller går på cricketmatcher vet vad en resultattavla är .
En resultattavla visar resultaten - den måste vara uppdaterad , tydlig och synlig .
Jag är övertygad om att kommissionär Vitorino kommer att se till att detta sker .
När de sex månaderna närmar sig sitt slut , hoppas jag att musiken fortfarande spelar och att de europeiska medborgarna fortfarande lyssnar .
Herr talman !
Jag vill välkomna rådets ordförande och hans kollega från justitiedepartementet , Costa , och tacka dem för det välkomnande de gav mitt utskott i Lissabon förra veckan och de konstruktiva sammanträden vi uppskattade .
Toppmötena i Amsterdam och Tammerfors har gett oss mycket arbete att utföra tillsammans , som det utmärkta resolutionsförslag som utarbetats av Terrón visar i dag .
Jag skulle vilja ta upp tre korta frågor .
Den första handlar om att vi behöver ett moget samtal mellan rådet och Europaparlamentet .
Det är knappt sex månader sedan det genom Amsterdamfördraget blev obligatoriskt för våra två organisationer att arbeta tillsammans ; vi har bedömt varandra , vi har haft några smågräl , men vi måste arbeta effektivt tillsammans .
Låt oss sluta med skuggboxningen .
Låt oss sluta med de omständliga charaderna och börja respektera de åtaganden som vi tagit på oss enligt fördragen och den tid det tar för en fullständigt demokratisk debatt .
Låt oss delta i era diskussioner om både politik och förfaranden .
Låt oss inte låtsas som om de nationella parlamenten kan utöva någon effektiv demokratisk kontroll över regeringsverksamheten inom detta område .
Min andra fråga handlar om att vi behöver en kommission som har tillgång till lämpliga resurser .
Vi har inrättat ett nytt generaldirektorat , ändå har detta bara 70 anställda .
Det finns ett avtal om att fördubbla denna siffra , men jag har förstått att inte en enda person har anställts ännu .
Vi ger kommissionen en tung uppgift , inte minst rörande utarbetandet av " resultattavlan " .
Rådet och parlamentet måste samarbeta för att tillhandahålla de resurser som kommissionen behöver .
Till sist , om debattinnehållet , välkomnar jag det faktum att ordförandeskapet placerat området för frihet , säkerhet och rättvisa högst upp på sin dagordning .
Alla goda ting äro tre , i synnerhet inom vårt politikområde .
För tvåhundra år sedan var det frihet , jämlikhet och broderskap och allt gick mycket bra ända tills olika vänsterregeringar satte jämlikheten över de andra .
Nu är det frihet , säkerhet och rättvisa och jag hoppas att de nuvarande vänsterregeringarna tar intryck av kommissionär Vitorinos ord och motstår frestelsen att sätta säkerheten - hur viktig den är - över de precis lika viktiga behoven i samband med frihet och rättvisa .
Kära kolleger !
Även om det är lämpligt att erinra om de viktigaste genomförandena i den europeiska uppbyggnaden av ett område för frihet , säkerhet och rättvisa , återstår fortfarande mycket att göra .
EG-domstolens roll är fortfarande alltför begränsad och överföringen till gemenskapsnivå förblir ofullständig .
Det räcker med att titta på Belgiens unilaterala beslut att återupprätta gränskontrollerna .
Beslutet att upprätta en stadga över de grundläggande friheterna är positivt , men det är svårt att förutse om dess innehåll och dess rättsliga omfattning , tvingande eller symbolisk , skall omfatta alla medborgare , oavsett nationalitet , eller utesluta vissa .
Man kan bara beklaga den totala avsaknaden av framsteg när det gäller det europeiska medborgarskapet och politiska rättigheter för alla invånare i Europa .
Även om handlingsplanen från högnivågruppen syftar till att i framtiden begränsa migrationsströmmen , förbättrar dessa planer inte på något sätt situationen för de mänskliga rättigheterna , de offentliga friheterna eller den ekonomiska situationen i de berörda länderna .
Vi vet att klausuler om återintagande finns i samarbets- och associeringsavtalen .
Men de utgör ett allvarligt hot mot principen om icke-avvisning .
Man måste också notera att dessa bestämmelser antagits inom rådet genom ett förfarande utan debatt och utan att parlamentet rådfrågats .
Det grundläggande problemet är ändå ....
( Talmannen avbröt talaren ) .
Herr talman !
Jag vill i likhet med mina kolleger välkomna rådets företrädare , såväl som kommissionsledamoten .
Jag tackar dem för deras uttalanden i kammaren .
I stället för att ta upp de redan diskuterade områdena , vill jag ta upp ett specifikt ämne : Narkotikafrågan och hur vi tar itu med den omfattande drogkulturen i våra samhällen .
Jag vänder mig särskilt till det portugisiska ordförandeskapet och uppmanar detta att bygga vidare på en del av det fantastiska arbete som utfördes av det finländska ordförandeskapet när det gällde att utarbeta samordnade planer och åtgärder mellan medlemsstaterna .
På den internationella sidan har vi redan börjat tillämpa planer för att bekämpa narkotikasmuggling , penningtvätt osv .
Men vi måste föra ned det på ett mer mänskligt plan : Att ge hjälp till de som försöker sluta med droger och ge dem lämpliga kontroller och lämpliga mekanismer för rehabilitering ; för det andra , att vidta samordnande åtgärder inom polisen och det rättsliga området vad gäller gemensamma straff och gemensam lagstiftning ; för det tredje , att genomföra en informations- och medvetandehöjande kampanj för yngre personer ; och en gång för alla stoppa användningen av de mycket farliga orden " normalisering " och " skademinskning " , och visa att all avmattning rörande vår beslutsamhet att se till att narkotika inte blir lagligt måste vara för medborgarnas bästa .
Herr talman !
Jag skulle vilja använda de futtiga sekunder talartid jag fått till att påpeka för kommissionens företrädare eller påminna honom om att regeringen i medlemsstaten Belgien just nu för en politik som innebär att tusentals och måhända tiotusentals illegala invandrare blir legaliserade , kommer att få permanent uppehållstillstånd , rätt till familjeåterförening , och så vidare .
Det är en åtgärd av den belgiska regeringen som är en flagrant överträdelse av Schengenavtalet .
Den 23 december lämnade jag in ett skriftligt klagomål om det till kommissionär Vitorino .
Jag skulle vilja be honom överväga det klagomålet och inom överskådlig tid tala om för mig vilka åtgärder kommissionen skall vidta för att straffa den belgiska statens överträdelse av Schengenavtalet enligt artikel 226 i avtalet .
Herr talman , mina värderade herrar från Portugal , särskilt rådets företrädare !
Ni befinner er i en situation där ni är ställda inför stora förväntningar från vår sida .
Jag vill med ett exempel visa hur ni rätt snabbt skulle kunna uppfylla dessa förväntningar , i vart fall inom ett begränsat segment .
Det handlar om Eurodac .
Ni minns att vi här i Europaparlamentet med stora förväntningar i december beslutade att Eurodac skall förverkligas som förordning och system , men också som instrument för gemenskapen ; detta behöver vi omgående för att få stopp på fenomenet med upprepade asylansökningar , för att få ett instrument mot laglösheten och framför allt för att klart kunna avgöra vilket medlemsland som bär ansvaret för ett asylförfarande .
Vi har klart tagit ställning för ett införande av detta instrument ; införandet kan ske via ett verkställande utskott som , tillsammans med motsvarande databas , bör vara knutet till kommissionen .
Vi var av åsikten att Eurodac borde förverkligas .
I Tammerfors var man av åsikten att Eurodac borde förverkligas .
Men redan vid nästa toppmöte i december valde rådet att ta ett steg tillbaka genom att besluta - vilket vi bestämt motsätter oss - att befogenheten att genomföra det skall ligga kvar hos rådet , att regelkommittén skall ligga hos rådet samt att Gibraltar om möjligt kan sättas in som ett påtryckningsmedel .
Detta är ett typexempel på hur arbetet inte bör ske .
Den enträgna begäran jag har för min partigrupps räkning är att ni gör allt som står i er makt för att omgående och snabbt förverkliga Eurodac som ett instrument för bekämpande av laglöshet och missbruk av asylreglerna samt som ett instrument för att åstadkomma snabba asylförfaranden .
Om ni i dag kunde säga oss hur ni tänkt gå tillväga skulle det vara mycket värdefullt för oss .
( Applåder ) Herr talman , herrar ministrar , herr kommissionär ! 1999 års skörd av beslut var verkligen riklig .
Så riklig , skulle jag vilja säga , att det blir svårt att ta hand om den , det vill säga att genomföra besluten .
Jag syftar särskilt på rådet och på medlemsstaternas slapphet att genomföra det som man bestämmer gemensamt .
Året som gick kännetecknades emellertid av flera positiva och avgörande beslut , till exempel trädde Amsterdamfördraget i kraft , Schengenavtalet införlivades i gemenskapspelaren , rådet beslutade i Köln att utarbeta en europeisk stadga för grundläggande rättigheter och vid det extra rådstoppmötet i Tammerfors förband sig medlemsstaterna att följa vissa gemensamma riktlinjer , prioriteringar och mål , med avsikten att skapa ett gemensamt område för frihet , säkerhet och rättvisa .
Samtidigt som vi erkänner de framsteg som har gjorts , betonar vi , som europeiskt parlament , den ovilja som har observerats hos rådet att genomföra besluten på många områden , bristen på samsyn och , framför allt , bristen på öppenhet och samarbete med Europaparlamentet .
Som jag sade märker ni kanske att Europaparlamentet inte är berett att spela endast observatörens roll .
Det kommer inte heller att upphöra med att ställa besvärliga frågor , som till exempel om hur långt ni är beredda att gå och vilka lagstiftningsåtgärder och andra åtgärder ni kommer att vidta för att bekämpa skammen med prostitution , barnpornografi på Internet , narkotikan och den organiserade brottsligheten .
Kommer ni att arbeta för en gemensam asyl- och invandringspolitik ?
Vad kommer ni att göra för att integrera invandrarna socialt , återförena familjer och ge tillgång till rättigheter och skyldigheter som är likvärdiga dem som gäller för medborgarna i unionen ?
Kanske kommer ni att bli tvungna att överge era traditionella konservativa åsikter om flyktingar och invandrare , inför den nya demografiska ordningen som beskrivs av FN : s sakkunniga .
Jag har stora förväntningar på det portugisiska ordförandeskapet .
Herr talman !
Jag välkomnar mycket , faktiskt det mesta , av vad som sagts under denna debatt .
Men jag vill att vi iakttar försiktighet .
Vi riskerar att få för många , inte för få , rättighetsstadgor i denna gemenskap : Konventioner på nationell , unions- och europeisk nivå ; det är inte får få domstolar som har det sista ordet om våra rättigheter , utan möjligen för många - vi har domstolen på andra sidan floden och domstolen i Luxemburg .
Det finns också domstolar i Karlsruhe , Lissabon , Dublin och Edinburgh .
Vi måste se till att det vi gör är förnuftigt .
Vi får inte skapa förvirring och konflikter när det gäller domsrätten i samband med rättigheter , för detta skulle vara skadligt för friheten , rättvisan och säkerheten .
Vi måste , kort sagt , ha och behålla högsta möjliga gemensamma standarder och hitta sätt att säkerställa dessa .
Men vi måste alltid ta hänsyn till subsidiaritetsprincipen .
Precis som alla andra i denna kammare vill jag ha frihet , säkerhet rättvisa .
Jag vill inte se att dessa värden degenererar och skapar övercentralisering , kaos och förvirring .
Fru talman , kära ledamöter !
Mycket snabbt skulle jag vilja säga följande : i ledamöternas inlägg har flera frågor ställts om det portugisiska ordförandeskapet .
Parlamentets talman fick oss att känna att den tid vi förfogar över är mycket kort och därför föreslår vi , jag och min kollega från justitiedepartementet , att vi objektivt besvarar alla frågor som ställs här , under mötet med det parlamentariska utskottet där vi kommer att närvara nästa vecka .
( Ihållande applåder ) Tack så mycket , herr minister !
Jag förklarar debatten avslutad .
Herr talman !
Jag tackar rådet för såväl det muntliga som det skriftlig svaret .
Effektiviteten är verkligen anmärkningsvärd .
Det ger mig några sekunder extra för jag ville föreslå rådet att vi fortsätter att debattera frågan nästa gång utskottet för medborgerliga fri- och rättigheter och inrikesfrågor träffas .
Då får vi tillfälle att kommentera de här svaren och uttala vår oro även inför kommissionen .
Personligen är jag glad för en del av svaren , som exempelvis de känsliga frågorna om Schengen eller Europolkonventionen , som vi hoppas kommer att revideras , och jag gläds över justitieministerns ord i den meningen att den skall försöka underställas den dömande maktens jurisdiktion .
Jag hoppas att man gör detsamma när det gäller den parlamentariska kontrollen Ärade företrädare från rådet , inom en månad kommer vi att lägga fram en resolution här i kammaren för votering .
Med det goda humör som ni har visat prov på i dag , så är jag säker på att det första som kommer att hända i det här nya klimatet av samförstånd är att ni kommer att beakta resolutionsförslaget .
 
Frågestund ( rådet ) Nästa punkt på föredragningslistan är frågor till rådet ( B5-0003 / 2000 ) .
Fråga nr 1 från ( H-0780 / 99 ) : Angående : Kärnkraftverk byggs på jordbävningsutsatta områden i Turkiet I Turkiet inträffade nyligen två jordskalv med en styrka på mer än magnitud 7 på Richterskalan .
Det är mycket oroande att Turkiet envetet tänker bygga några synnerligen kostsamma kärnkraftverk inom området Akkuyu samtidigt som energin från Atatürkdammarna exporteras till tredje land och EU ger ut pengar på att reparera de skador som uppstått vid jordbävningarna , i en situation där gemenskapen skär ner sin budget .
De turkiska kärnkraftsplanerna tar ingen hänsyn till de faror som kan uppstå för invånarna och ekosystemen i Turkiet och omgivande länder och de inger också misstankar om att Turkiets militära och politiska ledning på förhand utarbetat hemliga planer om att skaffa en teknik som skall bereda möjligheter till kärnvapenutveckling .
Det bör erinras att Turkiet söker bygga reaktorer som är av kanadensiskt ursprung och motsvarar de reaktorer som Indien och Pakistan anskaffat .
Vad tänker rådet göra för att kärnkatastrofer skall kunna undvikas och kärnvapenspridning förhindras till ett land som vill bli medlem av EU och som ger ut stora summor på kärnkraftsprogram men samtidigt tar emot ekonomiskt bistånd från EU ?
Herr talman !
Rådet vill klargöra att Turkiet har skrivit under konventionen om kärnsäkerhet , vars mål ligger i linje med den oro som uttrycktes av ledamoten .
Denna konvention , som trädde i kraft den 24 oktober 1996 , har just som syfte att uppnå en hög internationell kärnsäkerhet genom nationella åtgärder och genom internationellt samarbete , liksom att vid kärnkraftsanläggningarna etablera och upprätthålla ett skydd mot potentiella radiologiska risker för att skydda människor , samhälle och miljö mot skadlig joniserande strålning från denna typ av anläggningar .
Konventionen omfattar som bekant också skydd mot olyckor med radiologiska konsekvenser och ett minskande av dessa effekter när den här typen av olyckor inträffar .
Jag skulle dessutom vilja påpeka för ledamoten att Turkiet , som ansökarland till Europeiska unionen , förr eller senare , och detta är ett villkor innan anslutning - och jag tror att denna punkten är viktig - , i sin egen föranslutningsstrategi måste anta en politik som gör att landet i tid kan godta gemenskapslagstiftningen i helhet , inklusive alla bestämmelser som gäller för kärnsäkerhet .
Tack så mycket för svaret .
Jag skulle dock vilja tillägga följande .
Med denna enhet kommer Turkiet att öka sin energipotential med bara 2 procent .
Det sägs emellertid att Turkiet vill skaffa reaktorer av Candutyp , likadana som Pakistan och Indien har och med vars hjälp de har framställt kärnvapen .
Mot den bakgrunden måste saken undersökas , eftersom den känsliga situationen i Kaukasus kan leda in många i konstiga tankebanor .
För det andra , angående anläggningarnas säkerhet .
I regioner med stor jordbävningsfara räcker det inte med att vi har starka , jordbävningssäkra hus , för vid denna slags situationer - och jag säger er detta som ingenjör - använder vi modeller för att undersöka följderna av olika faror .
Vi kan emellertid inte göra modeller av kärnkraftsanläggningar i drift .
Det går inte .
Därför kan man a priori och på förhand säga att det inte går att ha kärnkraftsanläggningar i regioner med stor jordbävningsfara .
Av den anledningen , och eftersom Turkiet nu står på tröskeln till Europeiska unionen , måste vi hjälpa landet att bli ett säkerhetens , fredens och samarbetets land i regionen .
Det är vår roll , och det är målet med min fråga . - ( PT ) Herr talman !
Jag medger att de argument ledamoten framför är befogade .
Det handlar i verkligheten om en mycket känslig fråga .
Det är alltså en fråga , som ni förstår , som inte bara gäller Turkiet i sin närhet till den nuvarande Europeiska unionen , det gäller också andra stater som vi har förbindelser med genom vårt eget grannskap .
Vi förstår er oro och vi kommer att ta hänsyn till den , främst inom ramen för de framtida kontakterna med Turkiet när vi fastställer själva dagordningen för anslutningsstrategin för Turkiet .
Denna fråga hör till våra huvudangelägenheter och Europeiska kommissionen kommer med all säkerhet att beakta den .
Herr talman !
Jag tror , beträffande Newton Dunns fråga , att det är allmänt känt , även om det är värt att nämna det så att det kan noteras , att rådets generalsekretariat sedan 1996 utarbetar en månatlig sammanfattning av rådets lagstiftningsakter .
I denna sammanfattning medföljer , som bekant , eventuella förklaringar till akterna , med rösterna mot , nedlagda röster och röstförklaringar .
Från och med maj 1999 ( det gäller alltså perioden efter att Amsterdamfördraget trätt i kraft ) innehåller denna sammanfattning även de akter där rådet inte agerar som lagstiftare , utom vissa akter av begränsad omfattning , som besluten av processuell natur .
I detta fall kan sammanfattningen också inkludera röstresultatet om rådet så beslutar .
Dessutom offentliggör generalsekretariatet i sina pressmeddelanden efter varje möte med rådet , genom tillämpning av den interna förordningen från 1993 därefter ersatt av just rådets beslut av den 31 maj 1999 , eventuella omröstningsresultat och röstförklaringar där rådet agerar som lagstiftare , liksom i andra fall , genom ett ad hoc-beslut som rådet själv fattar .
Efter Amsterdamfördragets ikraftträdande och i de fall rådet agerar som lagstiftare - denna skillnad är viktig vad gäller ministerrådsmötenas funktion - , offentliggörs resultaten och röstförklaringarna , liksom förklaringar i akten , på ett systematiskt sätt .
Då bestämmelserna för offentliggörande är de samma för utarbetandet av de månatliga sammanfattningarna av rådets akter som för pressmeddelandena , är de eventuella omröstningar som finns med i den ena eller den andra informationen precis samma , frånsett eventuella misstag som kan uppstå .
När det gäller Frahms och Sjöstedts frågor kan jag säga att de allmänna principer och begränsningar , enligt artikel 255.2 i fördraget med de ändringar som infördes genom Amsterdamfördraget , som för allmänhetens eller de privata intressenas skull måste reglera rätten att ta del av dokumenten , kommer att fastställas av rådet , som behandlar dem i en medbeslutandeprocess med detta parlament , utifrån ett förslag av Europeiska kommissionen , ett förslag som skall läggas fram - som ni känner till inom ramen för Amsterdamfördraget - inom en tidsfrist om två år efter Amsterdamfördragets ikraftträdande , det vill säga före 1 maj 2001 .
Eftersom rådet hittills inte har fått något förslag från kommissionen i denna fråga , förstår ni säkert att jag inte kan svara på de detaljfrågor som ledamöterna har tagit upp .
Tack , herr talman och tack , herr rådsordförande !
Jag är säker på att rådsordföranden är en mycket trevlig man och att han är mycket vänlig mot sin fru , sina barn och sin hund .
Ni måste emellertid förlåta mig om jag är litet skeptisk rörande det svar ni just gett mig .
Jag tror inte att de uttalanden som görs i rådet och omröstningsresultaten omedelbart finns tillgängliga för allmänheten .
Kan ni därför , före nästa sammanträdesperiod i februari , skriva till mig och berätta var jag kan hitta denna information på allmänhetens vägnar så snart som rådet har antagit lagstiftning , i stället för att vänta på att den skall offentliggöras veckor senare som pressmeddelande .
Kan ni skicka nämnda information till mig före nästa sammanträdesperiod ? - ( PT ) Herr ledamot !
Jag vill först säga att jag undanber mig personliga kommentarer av det slag som ni inledde er andra fråga med och om ni kan bespara oss dessa i framtiden skulle jag vara tacksam .
I det ni framförde ger ni oss idén att kritiken mot rådet , förutom att den är formulerad på ett mycket speciellt sätt vilket vi också noterar , inte handlar så mycket om ogenomskinligheten , om vi kallar den så , i lagstiftningsprocessen , utan snarare om en överdriven öppenhet .
Men jag skulle vilja säga , herr ledamot , att vi anser att resultaten av denna typ av arbete för öppenhet är klara och tydliga .
Vi tvekar inte , herr ledamot , att upprepa denna information skriftligt , men vi kan inte gå längre än vad vi säger eftersom det vi säger är precis det fördraget kräver .
Vi anser alltså att alla de element som rådets generalsekretariat förser allmänheten med är de viktiga element som krävs för att rådet skall fungera som lagstiftande myndighet .
Jag anser att rådet inte försökte svara på min fråga .
Jag frågade inte vad rådet ansåg om det förslag som kommissionen ännu inte har lagt fram , utan min fråga gäller den principiella tolkningen av artikel 255 i Amsterdamfördraget .
Medger den att man lagstiftar också om nationell öppenhetslag , inte bara om de tre institutioner i Europeiska unionen som anges där ?
Jag skulle gärna vilja ha ett svar på denna fråga .
Anser rådet att man på grundval av artikel 255 i fördraget kan reglera nationell öppenhetslagstiftning , dvs. inte den som avser EU : s institutioner ? - ( PT ) Herr talman !
Det svar ni fick var det svar som var möjligt att ge .
Jag vill emellertid säga följande : tolkningen av artikel 255 i fördraget är en tolkning som också måste vara knuten till subsidiaritetsprincipen .
Det finns för närvarande inget konkret förslag som gör det möjligt att arbeta med förordningen för denna artikel , och utan detta förslag är det inte möjligt att göra framsteg i frågan .
Hur som helst , den första tolkning vi gör är att artikel 255 inte gör det möjligt att arbeta på ett sätt som påverkar subsidiaritetsprincipen .
Jag är absorberad av det sätt på vilket rådet kämpar för de principer som finns i Amsterdamfördraget , och som handlar om att se till att medborgarna får en bättre möjlighet att delta i beslutsprocessen .
Hur gör man det när man samtidigt enligt kommissionens uttalande - det har läckt ut , så det är allmänt känt - säger att de anställdas tankefrihet sätts framför öppenheten , så att man inte kan få tillgång till arbetsdokument , rapporter , förslag osv . ?
Anser inte rådets företrädare att detta försvårar ett deltagande i den demokratiska beslutsprocessen ?
Fru ledamot !
Den fråga ni har ställt är av största vikt och vi diskuterade den länge under senaste regeringskonferensen .
Och jag vill säga er en sak : gemenskapsinstitutionernas öppenhet fungerar inte bara " utåt " , de fungerar också " mellan " gemenskapens institutioner .
Det vill säga , det finns saker i formen och arbetsprocessen i gemenskapsinstitutionerna som inte är tillgängliga för andra institutioner , och det gäller inte bara mellan kommissionen och parlamentet , det gäller också mellan kommissionen och rådet .
Detta ämne har alltså redan tagits upp och diskuterats flera gånger .
Europaparlamentet kommer att ha möjlighet att medverka i den grupp som förbereder nästa regeringskonferens .
Det är en öppen fråga .
Utformningen av och den reella öppenheten i de europeiska institutionernas verksamhet är en fråga av största betydelse och det är en fråga som , enligt min mening måste analyseras än en gång , främst inom ramen för nästa regeringskonferens , detta är vi helt på det klara med , och vi menar att de ledamöter som deltar i denna förberedande grupp , får ännu ett tillfälle att ta upp denna fråga .
Jag tycker att kommissionens förslag bör innehålla element för att skapa en större öppenhet i förhållande till verksamheten i de olika institutionerna , men jag menar att det alltid finns utrymme för förbättringar i denna fråga .
För vår del är vi beredda att behandla de förslag som läggs fram på detta område .
Det är en väldigt viktig fråga som Jonas Sjöstedt och andra har ställt .
Vi har en offentlighetsprincip i Sverige som stärker demokratin och som ser till att det blir en bra dialog mellan medborgare , beslutsfattare och myndigheter .
Vi är väldigt måna om att även EU skall gå åt detta håll , och det står även i Amsterdamfördraget .
Parlamentet antog ett betänkande av Lööw för ett eller ett par år sedan som är väldigt viktigt i detta sammanhang .
Däri varnades det för att den kommande processen skulle leda till inskränkningar i medlemsländernas offentlighet .
Nu kan vi se att det kanske finns ett visst fog för denna varning från parlamentet .
Jag vill fråga rådet om rådet har förståelse för denna varning , med tanke på det som vi nu har sett i arbetsdokumenten från kommissionen . - ( PT ) Fru ledamot !
Vi bör alla vara medvetna om en sak : mellan rådet och parlamentet , mellan rådets medlemmar och medlemmarna i detta parlament råder det inte nödvändigtvis någon klyfta vad gäller fördelarna eller nackdelarna med öppenheten .
Ibland skapar man sig en idé om att rådet är ett högkvarter för slutenhet och parlamentet är ett högkvarter för öppenhet .
Det är inte sant .
Vi är lika angelägna som ledamoten om institutionernas sätt att fungera och vilken effekt detta funktionssätt har utåt .
Vi delar alltså samma oro och tolkar principerna på samma sätt .
Det som kan hända , fru ledamot , är att vi på sina håll inte har samma tolkning på hur arbetet med öppenheten exakt skall gå till i förhållande till en verklig öppenhet .
Det vill säga , ofta är tanken att spridningen av en viss typ av dokument , och att ett öppet sätt att arbeta i vissa institutioner är en faktor som fungerar till förmån för demokratiseringen av dessa institutioner , en farlig tanke eftersom detta ofta inte sker .
Vi vet - och jag vill inte breda ut mig för mycket om det - , vi vet att vi , när öppenheten ibland går över vissa gränser , hamnar i en situation där samtalen och förhandlingarna sker i korridorerna .
Det finns en allmän balans i frågan om öppenhet .
Och det finns en balans som går precis mellan realism och demagogi .
Jag lyssnade med stor uppmärksamhet till det som Seixas da Costa sade om öppenheten och regeringskonferensen .
Min fråga är om jag av det som Seixas da Costa sade , de intressanta sakerna om öppenheten och regeringskonferensen , kan dra slutsatsen att det portugisiska ordförandeskapet förbinder sig att arbeta och kämpa för en utvidgning av regeringskonferensens dagordning .
För undersökningen av frågan om " öppenhet " med avseende på institutionernas funktion kan hur som helst inte gömmas undan på något ställe och i några frågor eller i några korridorer - även om också jag inser korridorernas betydelse .
Den kräver en särskilt punkt på regeringskonferensens dagordning , vilket innebär en utvidgning av denna . - ( PT ) Herr talman !
Frågan om öppenhet är en fråga som naturligtvis har att göra med institutionerna .
Denna regeringskonferens sätter i gång med en inriktning , åtminstone inledningsvis , på att få institutionerna att fungera bättre , särskilt med hänsyn till den önskan vi alla har om att de skall bli just mer demokratiska , öppna och effektiva .
Allt detta befinner sig dock inom en allmän ram , den allmänna ramen om en gemensam acceptans av alla lösningar vi kan finna för att genomföra dessa tre önskningar .
Det är uppenbart att denna öppenhet ständigt kommer att finnas med på den europeiska dagordningen och den kommer givetvis att vara med på denna regeringskonferens .
Det är en fråga som det portugisiska ordförandeskapet , det kan jag försäkra er , kommer att tas upp med medlemsstaterna och företrädarna för den grupp som förbereder konferensen .
Ordförandeskap bör i detta få stöd av Europaparlamentets ledamöter , vilka säkerligen är beredda att stödja detta förslag .
Därefter får vi se vilket resultat vi kan uppnå på ministernivå .
Vi bör dock tänka på att vi just har avslutat ett Amsterdamfördrag som godkändes i maj förra året , och att det där finns en mängd åtgärder för öppenhet som skall genomföras och som är på gång , och frågan är om det är för tidigt att sätta i gång ett nytt arbete om öppenhet .
Jag tycker trots allt att detta är en fråga som alltid bör vara med på dagordningen , eftersom det finns en viss märkbar sensibilitet hos allmänheten angående detta , och för att det i verkligheten handlar om behovet att göra de europeiska institutionernas organ ansvariga inför medborgarna .
För vår del kommer den att finnas med .
Vi får se om vi uppnår enhällighet för detta .
Fråga nr 5 från ( H-0785 / 99 ) Angående : Förslag till förordning som anger total tillåten fångstmängd för vissa fiskarter ( i detta fall ansjovis ) för år 2000 Enligt de senaste rapporterna från Internationella havsforskningsrådet ( ICES ) är den aktuella situationen i ICES-zon VIII kritisk för ansjovisbestånden .
Har rådet ( fiske ) och kommissionen undersökt hur ansjovisbestånden i zon VIII har påverkats av att ICES-zonerna IX och X och CECAF : s ( fiskerikommittén för östra centralatlanten ) zon 34.1.1 överlåtits från Portugal till Frankrike ( fiskekvoterna överskrids med 5 000 ton / år ) ?
Har man undersökt Frankrikes ansvar för den nuvarande situationen och för möjliga framtida ekonomiska och sociala konsekvenser för fiskesektorn ?
Anser rådet att det är godtagbart att tillåta fortsatt överfiske som strider mot den ursprungligen fastställda totalt tillåtna fångstmängden på 33 000 ton / år , när det råder en så kritisk situation för ansjovisbestånden ?
När tänker rådet vidta några åtgärder , och vilka kommer dessa att vara , för att behandla det kritiska läge som råder för ansjovisbestånden och sätta det i samband med överlåtandet av de portugisiska kvoterna och med principen om relativ stabilitet ?
Herr talman !
Det portugisiska ordförandeskapet har allt intresse av att besvara denna fråga på ett fullständigt sätt , eftersom det också handlar om ett problem som berör Portugal på ett positivt sätt , och jag skall förklara hur .
Rådet är medvetet om den kritiska situationen för ansjovisbestånden i havet utanför Kantabrien som ledamoten tar upp .
Ändå ansåg de medlemsstater som utför detta fiske , det vill säga Frankrike , Spanien och Portugal , vid det senaste rådsmötet ( fiske ) förra året , den 16 och 17 december , att tillämpningen av försiktighetsprincipen som fastställer en minskad tillåten totalfångst från 5 000 ton till 2 000 på förslag av kommissionen , var överdrivet försiktig .
Man kom då fram till en kompromisslösning för att nå en balans mellan behovet att minska de biologiska riskerna , alltså påverkan på fiskbestånden , och de socioekonomiska svårigheterna som orsakas av ett begränsat fiske , med en fastställd tillåten totalfångst på en mellannivå om 16 000 ton i stället för 33 000 som var förutsett för 1999 .
En revidering planerades också i ljuset av ny information av vetenskaplig karaktär angående bevarande av arterna som man hoppas skall bli klar under första halvåret i år .
För det södra ansjovisbeståndet , i ICES-zonen IX , fastställdes den tillåtna totalfångsten till 10 000 ton för år 2000 mot 13 000 ton för 1999 .
Förändringarna av fiskemöjligheter mellan Portugal och Frankrike minskades proportionellt från 5 008 ton för 1999 till 3 000 ton år 2000 , i de franska fiskevattnen .
Jag skulle vilja nämna att denna överföring inte kommer att öka fisketrycket på ansjovisbeståndet i sin helhet , inom hela gemenskapens fiskeområde .
Och i enlighet med principen om relativ stabilitet , tilldelades Spanien 90 procent av beståndet och Frankrike bara 10 procent av fördelningsnyckeln för ansjovisfisket i havet utanför Kantabrien .
Utan en överföring till de portugisiska fiskevattnen , skulle den tillåtna totalfångsten i havet utanför Kantabrien behöva ökas tio gånger för att ge Frankrike ett adekvat fiske .
Detta är skälet till att jag anser att det finns ett positivt element i Portugals fall .
Det är uppenbart att denna lösning skulle skada fiskbeståndet ännu mer än den risk ledamoten talade om , men vi förstår det .
Herr rådsordförande !
Jag måste säga att ert uttalande ingalunda har lämnat mig tillfreds .
Jag förstår att Portugal berörs av detta .
Det är enligt min mening som ett attentat mot det sunda förnuftet och intelligensen att 80 procent av den ansjovis som fiskades i portugisiskt vatten efter avtalet mellan medlemslandet Portugal och Frankrike i stället börjar fiskas i Biscayagolfen och att ministerrådet vidhåller att detta varken påverkar ansjovisbeståndet där eller i Biscayabukten .
Allt sedan 1995 har vi visat att den här omflyttningen är rena galenskapen och om Portugal och Frankrike vill träffa en överenskommelse så får de väl det , men ansjovisen skall fångas i portugisiskt vatten och inte i Biscayagolfen .
I dag visar vetenskapliga studier att ansjovisbestånden i Biscayagolfen är utrotningshotade .
Och nu kommer inskränkningar i de ansjoviskvoter som skall gälla för Biscayagolfen .
Ärade rådsministrar , jag vet inte om ni är medvetna om att ni har ett ansvar för det som hänt under de här åren men också för år 2000 när det gäller de tusentals familjer på norra delen av iberiska halvön som lever av ansjovisfiske . - ( PT ) Jag skulle vilja säga , herr ledamot , att EG-domstolen i sin dom den 5 oktober 1999 , beslutade att denna överföring , en överföring som godkändes , var i överensstämmelse med de principer som fastslås i rådets förordning 37 / 60 / 92 och främst artikel 9.1 vilken säger att medlemsstaterna kan byta hela eller delar av sina tilldelade fiskerättigheter .
Domstolen uttalade också att principen om relativ stabilitet inte hade kränkts eftersom ansjoviskvoten som tilldelats Spanien i underkategori 8 behölls på 90 procent och Frankrikes kvot på 10 procent .
Dessutom , herr ledamot , är domstolen av den åsikten att överföringen mellan Portugal och Frankrike inte kränker principen om rationellt och ansvarsfullt fiske i hav och levande vattendrag eftersom fisketrycket i underkategori 8 och 9 inte ökar eller innebär någon negativ påverkan för den allmänna kvoten av de resurser som tilldelats Spanien .
I enlighet med detta , herr ledamot , upprepar rådet sin åsikt att utan denna överföring , skulle en hänsyn till Frankrikes fiskemöjligheter göra att ansjovisfisket i Biscayabukten öka .
Rådet upprepar alltså , herr ledamot , sin åsikt om att fisketrycket skulle vara större och mer skadligt för fiskbestånden än den lösning som nu har valts .
Konkret utgör 3 000 ton 57,5 procent av Portugals fiskemöjligheter under 2000 , mot 5 008 ton , eller 73,9 procent 1999 .
Dessa siffror utgör , enligt vår åsikt och rådets perspektiv , en verklig förbättring vad gäller bevarande jämfört med en nivå på 80 procent som fastställdes i rådets förordning 685 / 95 .
Fråga nr 6 från ( H-0788 / 99 ) : Angående : Åtgärder mot den fortgående etniska rensningen av Kosovos serber och romer Natos försvarsministermöte sände den 2 december 1999 ut en kraftfull appell genom vilken man kräver ett slut på den etniska rensningen av Kosovos minoriteter .
Europaparlamentet fördömer också i en av sina resolutioner , med hänvisning till de fruktansvärda våldshandlingar som riktats mot serber och romer , det fortsatta våldet mot den serbiska befolkningen och uppmanar de albanska ledarna i Kosovo att till fullo respektera FN : s beslut nr 1244 .
I denna resolution betonar parlamentet att de tidigare förföljelserna av albaner inte kan accepteras som ursäkt för " fortsatt dödande , kidnappningar , interneringar , maktmissbruk , trakasserier , hotelser , mordbränder , plundring , förstörelse av egendom och husövertaganden " etc .
Ämnar rådet - mot bakgrund av ovanstående B ta upp frågan om finansieringen av återuppbyggnadsarbetena i Kosovo till ny granskning , i enlighet med Europaparlamentets krav ?
Vilka övriga konkreta åtgärder ämnar rådet vidta för att få ett slut på den etniska rensningen ?
Herr ledamot !
Jag skulle vilja säga att jag har mycket sympati för den oro som ligger bakom er fråga .
Vi delar verkligen den oro ledamoten hyser inför den hotfulla situation som råder i Kosovo för de etniska minoriteterna , både den serbiska befolkningen och romerna , och som handlar om fortsatt diskriminering , förföljelser och hot på detta territorium .
Rådet betonar alltid att det är nödvändigt att döma de som har begått och de som fortsätter att begå sådana handlingar Rådet upprepade också , i sina slutsatser från december , att det var nödvändigt med en fullständig tillämpning av säkerhetsrådets resolution 12 / 99 och har systematiskt stött Bernard Kouchners arbete för att införa åtgärder som kan garantera ett effektivt skydd för minoriteterna i området , och särskilt en effektiv tillämpning av åtgärder som gör det möjligt att bevara det multietniska samhället i området .
I de kontakter vi har haft med de mest framstående politiska företrädarna för Kosovos albaner , och dessa kontakter togs alldeles nyligen av den portugisiske premiärministern , har vi framhållit att förföljelserna av den serbiska befolkningen , den zigenska befolkningen och andra etniska grupper är fullkomligt oacceptabel .
Detta kommer inte att tolereras och det bör genast upphöra .
Detta meddelades tydligt och upprepade gånger till Kosovos ledares att det internationella stödet till stor del är avhängigt av behandlingen av de icke-albanska etniska minoriteterna .
Jag anser att denna punkt är av största vikt , denna känsla av förutsättning som ligger i Europeiska unionens ståndpunkt kommer att vidmakthållas av rådet .
Vi har stött FN-uppdragets och den internationella säkerhetsstyrkans arbete i Kosovo för att förhindra nya våldsuttryck mot minoriteterna och att skydda de hotade befolkningsgrupperna .
Kafor och polisen Minuc ser som en av sina viktigaste uppgifter att på alla sätt få bort kränkningarna på grund av etniskt ursprung .
I detta sammanhang gläds rådet i sina slutsatser från december , åt det substantiella bidrag som Europeiska kommissionen har meddelat att den skall ge indirekt till normaliseringen av situationen tillsammans med liknande bidrag från medlemsstaterna .
Emellertid , herr ledamot , är rådet också medvetet om att alla medel som ges till internationellt ansvariga strukturer i Kosovo inte motsvarar de som vore önskvärda , när det gäller mobilisering i de olika medlemsstaterna , och detta begränsar den effektiva handlingsförmågan när det gäller dessa strukturer .
Vi kommer emellertid att koncentrera all vår uppmärksamhet på detta problem eftersom all trovärdighet för de albanska myndigheterna och strukturerna i området också beror på dessa strukturers förmåga att visa att de kan vidta åtgärder som garanterar ett multietniskt samhälle i området .
Jag skulle vilja tacka rådsordföranden .
Min åsikt - och allas vår åsikt , tror jag - är att Portugal , landets förre president , Soares , och landets regering intog en förnuftig och moderat hållning under bombningarna på Balkan .
Och dagens politiska uttalande om denna fråga är mycket positivt .
Det vill jag betona och välkomna .
Trots detta finns det anledning till oro , för samtidigt som det från Europeiska unionens sida finns goda och uppriktiga föresatser , är resultaten mycket små .
Den senaste tiden har vi tyvärr sett en utplåning av alla minoriteter - av serber , romer , turkar , kroater - i Kosovo , och vi frågar oss vad som kommer att hända .
Förenta nationernas och Kouchners uppdrag i Kosovo är ett misslyckande .
Det faktum att vi efter ett fullständigt krig som startades för att förhindra etnisk rensning nu förekommer etnisk rensning från den motsatta sidan är ett misslyckande .
Av den anledningen upprepar jag min fråga , om rådet har för avsikt att vidta mer konkreta praktiska åtgärder för att diskutera dessa frågor med Kouchner , som har ett mycket stort ansvar för den situation som i dag råder i Kosovo . - ( PT ) Herr Alavanos !
Jag kan inte hålla med er om det ni säger i den sista meningen om Kouchners ansvar , och jag skulle vilja urskilja två mycket viktiga nivåer : den struktur som införts i Kosovo är en struktur under FN : s beskydd .
Det är en struktur som Europeiska unionen har gett det stöd som varit möjligt och till vilket länderna i Europeiska unionen har bidragit på olika sätt .
Men det finns en sak vi inte kan förneka , det är att Kouchners ansträngningar för en normalisering av situationen i Kosovo är oerhört positiva ansträngningar .
Oberoende av om ledamoten kan tycka , vilket vi också gör , att vissa av resultaten , av skäl som inte haft att göra med Kouchner , av dessa ansträngningar inte har varit så effektiva som vi alla hade önskat .
Här måste vi göra en sista distinktion i ansvarsfrågan för Europeiska unionen och i detta fall främst mellan rådets möjliga handlingsförmåga i detta sammanhang , och det internationella samfundets ansvar , vilket har det allmänna ansvaret för situationen i Kosovo .
Europeiska unionens ansvar hör alltså till ett visst bestämt sammanhang .
Det är internationella samfundet , nämligen FN , som skall avkrävas ansvar för genomförandet av resolution 12 / 99 och särskilt för logiken i denna resolution och förenligheten mellan resolutionen och verkligheten .
Detta är frågor vi alla bör ställa oss , men det rätta forumet för dessa frågor är FN .
Herr talman !
Herr rådsordförande , jag välkomnar varmt era ord att ni har för avsikt att förbättra organisationen och att det handlar om att öka myndigheternas trovärdighet .
Jag tror att vi då också bör fundera över hur vi på bästa sätt skall presentera det för allmänheten .
Jag frågar mig därför : Finns det egentligen några idéer om hur vi kan bearbeta medierna på detta område , hur vi kan ge journalister utbildning och hur vi på ett bättre sätt kan informera allmänheten om fredlig samlevnad ?
Vi har försökt att ge materiellt stöd .
Vi har också försökt att på militär väg åstadkomma fred .
Hur ligger det till med våra strävanden att också arbeta med psykologiska omständigheter i detta krisområde och på så sätt ge bästa möjliga stöd ? - ( PT ) Herr ledamot !
Som jag sade förstår jag er oro .
Jag anser att det just nu och särskilt de senaste månaderna har skett en viss positiv utveckling vad gäller de medel Kouchner kan förfoga över för ett effektivt arbete .
Jag minns att jag hörde Kouchner under ett ministermöte med Europeiska rådet i denna fråga och många angelägenheter han då påtalade angående bristande medel för att lyckas övervinna vissa problem är i dag lösta , det vill säga , han har nu fått dessa medel .
Vi har framför allt två viktiga frågor : för det första , en ökad polisens resurser , vilket var en viktig fråga för att skydda civilbefolkningen , och särskilt vissa befolkningar , och ökade anslag för att främst kunna behålla vissa viktiga administrativa och operativa funktioner i processen .
Frågan , herr ledamot , och det är en fråga som vi alla borde ställa , och jag gjorde det nyligen på ett diplomatiskt sätt , gäller själva karaktären på säkerhetsrådets resolution 12 / 99 .
Jag vet att det är en mycket känslig fråga men vi är alla rädda att ifrågasätta den inneboende logiken i denna resolution och möjligheten att genomföra den .
Vi stöder helt och hållet dess fullständiga genomförande : Vi måste dock granska denna resolution - och troligen måste FN : s säkerhetsråd förr eller senare göra detta - , för att kunna bedöma , så som har skett i andra internationella strategiska scenarier , om en viss typ av agerande och en viss typ av omständighet och balans - alltså de omständigheter och balanser som ledde till att resolutionen antogs - , skall bibehållas eller ej i framtiden .
Vi bör , och detta sker från Europeiska unionens sida , se till att Kouchner får alla resurser , och ledamoten har rätt , vi måste regelbundet och öppet förklara för våra medborgare huruvida dessa resurser används på ett bra sätt eller ej .
Rådet tänker givetvis under det portugisiska ordförandeskapet komma med information i denna fråga .
Herr rådsordförande !
Jag är helt överens med er .
Problemet är inte herr Kouchner , utan den rättsliga grunden han arbetar utifrån , nämligen resolution 1244 .
Jag tror därför att det är unionens ansvar , dvs. ert , men också vårt , att börja arbeta för att komma förbi den provisoriska karaktären i resolution 1244 och tänka oss ett framtida scenario för hela regionen .
Jag tror att det är denna brist på definition av scenariot som åstadkommer eller gynnar de översvämningar , olyckor och mord som Alavanos talat om .
Avser rådet att ställa frågan om Kosovos definitiva status ?
Och om så är fallet , avser man att göra det i en allmän omdefiniering av regionen , och genom att så långt det är möjligt undvika att öka mikrostaterna , såsom vissa har tendens att göra , och genom att på nytt ena parterna , i detta fall Kosovo och Albanien ? - ( PT ) Det är uppenbart , herr ledamot , att rådet inte kommer att försöka förändra statusen för Kosovo utanför den ram som slås fast i säkerhetsrådets resolution 1244 / 99 .
Jag skulle vilja säga att hanteringen av denna fråga i säkerhetsrådet även väcker en annan ganska intressant fråga , den om hur Europeiska unionen skall företrädas i detta råd , och alltså huruvida Europeiska unionens representation i säkerhetsrådet följer bestämmelserna för den gemensamma utrikes- och säkerhetspolitiken eller inte .
Men detta skulle troligen ta mer än ett sammanträde med parlamentet för att diskutera .
Jag vill dock säga att vi anser att situationen i Kosovo är en situation som också handlar mycket om situationen i alla de länder och områden som omger Kosovo .
Situationen i Kosovo är en situation som inte kan lösas i sig , den måste lösas genom en allmän stabilitet i hela regionen .
Detta skall naturligtvis ske genom de åtgärder som vidtas inom ramen för Europeiska unionen , både för en stabilisering av situationen i Bosnien och Hercegovina , liksom för de nya förbindelser vi försöker skapa i form av avtal med Före detta jugoslaviska republiken Makedonien , samt även alla åtgärder av positiv karaktär som vi försöker genomföra i Albanien , och naturligtvis det tryck vi sätter på de serbiska myndigheterna främst genom stödet i projektet " Energi för demokratin " , som vi ger de serbiska kommuner med demokratiska strukturer .
Detta är de åtgärder som , i sin helhet och genom synergism , också kan leda till en anda som kan lösa situationen i Kosovo .
Situationen i Kosovo kan inte lösas om det inte finns ett allmänt stabiliseringsprojekt i regionen .
Eftersom frågeställaren är frånvarande , bortfaller fråga nr 7 .
Fråga nr 8 från ( H-0796 / 99 ) : Angående : Nytt INTERREG-initiativ Enligt kommissionens meddelande om INTERREG , om främjande av utveckling i städer , på landsbygden och längs kusterna , bilaga 2 punkt 1 , skall man tillåta renovering och utveckling av historiska stadscentrum med hjälp av gränsöverskridande åtgärder .
Däremot framgår det tydligt att bostäder inte skall omfattas .
På landsbygden finns det många bostäder som är av historiskt intresse , exempelvis små stugor , och man bör av flera skäl bibehålla landsbygdsbefolkningarna och locka folk att bo i landsbygdsområdena .
Håller inte rådet med om att dessa målsättningar därför skulle kunna understödjas genom att finansiera bostadsprojekt inom ramen för INTERREG ? , rådet .
( PT ) Herr talman !
Rådet , och jag skulle särskilt vilja säga det portugisiska ordförandeskapet , är oerhört medvetet om betydelsen av de problem som ledamoten fokuserar i sin fråga och jag vill säga att vi hela tiden ägnar all uppmärksamhet åt den gemensamma politiken för utveckling av landsbygden .
I detta sammanhang skulle jag vilja framhäva antagandet i maj 1999 , av ett nytt system för stöd till landsbygdens utveckling , vilket utgjorde gemenskapens referensram för en hållbar utveckling av landsbygden och det var , som ni vet , ett av de projekten inom ramen för förhandlingarna om agenda 2000 och i utvecklingen av jordbruksfrågornas hantering på gemenskapsnivå .
Genom Europeiska utvecklings- och garantifonden för jordbruket ( EUGFJ ) , är denna gemenskapens stödram inriktad på stöd till att vända tendensen till utbredning av ödemark vilket ledamoten helt befogat tar upp i sin fråga .
Även Europeiska investeringsfonden ( EIF ) , bidrar till detta arbete med att främja den ekonomiska och sociala sammanhållningen genom att rätta till de största regionala ojämlikheterna och delta i utvecklingen och omställningen av landsbygden .
Det är lämpligt att tänka på att EIF har bidragit på samma sätt till främjandet av en hållbar utveckling av landsbygden som att skapa hållbar sysselsättning .
Det är dessa gemenskapsinstrument i sin helhet som gör det möjligt att arbeta i en politik för landsbygdsutveckling som i dag är ett utvecklingsområde och en inriktning i den gemensamma jordbrukspolitiken å ena sidan och regionalpolitiken å den andra .
Vi anser att detta , inom begreppet mångsidighet som i dag är knutet till utvecklingen av den gemensamma jordbrukspolitiken , är en av de grundläggande frågorna och EUGFJ : s garantisektion spelar naturligtvis här en fundamental roll .
Fråga nr 9 från ( H-0798 / 99 ) : Angående : Jordbruk och ordförandelandet Portugal Kan rådet ange ordförandelandet Portugals prioriteringar för den gemensamma jordbrukspolitiken för det närmaste halvåret och de åtgärder det anser vara nödvändiga för att öka konsumenternas förtroende för jordbrukssektorn och jordbruksprodukter , efter att detta förtroende har minskat på grund av den senaste tidens hälsorelaterade farhågor ? , rådet .
( PT ) Frågan som ledamoten ställer om den gemensamma jordbrukspolitiken är en fråga som berör oss nära , och det är värt att alltid ha den med i diskussionerna i denna kammare , för vi kommer troligen att ha mycket att diskutera i detta ämne i framtiden .
Under det portugisiska ordförandeskapet måste vi fortsätta debattera arbetet med den gemensamma jordbrukspolitiken , genom att anta några av de gemensamma organisationerna av marknaden med hänsyn till en harmonisk utveckling av unionens landsbygdsområden och en garanti om en positiv utveckling av jordbrukarnas inkomster , med särskild uppmärksamhet på de åtgärder som kan få följder för de små familjejordbruken .
Det portugisiska ordförandeskapet kommer naturligtvis också , om den nya rundan i Världshandelsorganisationen inleds under dess ordförandeskap , en sak som är långt ifrån säker , att försäkra sig om att befästa närvaron av gemenskapsproduktionen på de internationella marknaderna och en bättre balans mellan gemenskapens jordbruksprodukter som exporteras , samt bevarandet av ett mångsidigt europeisk jordbruk , vilket jag redan har nämnt .
Det portugisiska ordförandeskapet kommer också att lägga vikt vid en fördjupning av politiken för livsmedelssäkerhet och detta tog den portugisiske utrikesministern och rådsordföranden för Europeiska unionen , upp i dag på förmiddagen .
Vi anser att livsmedelssäkerhetens roll , framför allt när det gäller folkhälsan , är en mycket viktig sak som vårt ordförandeskap skall arbeta med , det utgör för övrigt en av prioriteringarna i vårt program .
Vi kommer att arbeta med detta inom fyra parallella områden inom ramen för Agrifin-rådet , rådet ( hälso- och sjukvård ) , rådet ( konsumentfrågor ) och rådet ( inre marknaden ) .
Det portugisiska ordförandeskapet kommer i juni i år , under Europeiska rådet i Santa Maria da Feira , också att lägga fram en rapport på detta tema , framför allt i ljuset av det som kommissionen för några dagar sedan presenterade i sin vitbok .
Vi tycker att det arbete vi skall göra från och med nu för att konstituera en europeisk byrå är ett viktigt arbete för att skapa trovärdighet för den inre marknaden och för att stabilisera det egna förtroendet inom denna marknad , upplösa vissa spänningar mellan medlemsstater på detta område och till och med , varför inte säga det rakt ut , att skapa en gemensam hållning från Europeiska unionens sida i sina förbindelser med tredje land på områden som handlar om livsmedelssäkerhet .
Detta är det arbete vi skall försöka genomföra under det portugisiska ordförandeskapet och vi hoppas i slutet kunna presentera resultatet av detta arbete .
Jag vill tacka rådets ordförande för hans svar .
Jag är säker på att han är medveten om det mycket allvarliga hotet mot den europeiska modellen , som grundas på familjejordbruk , i huvudsak mot de jordbrukare som sysslar med nötkötts- och fårköttsproduktion och som nu förväntas sälja sin produktion till eller under produktionskostnad .
Jag vill fråga vilka nya åtgärder som rådet kan vidta för att skydda deras intressen under de kommande samtalen inom Världshandelsorganisationen , i synnerhet mot den stordrifts- och industriliknande produktion som sker i Förenta staterna och Nya Zeeland där stordriftsfördelarna gör det oerhört svårt för de europeiska jordbrukarna att skapa konkurrenskraftiga familjejordbruk och där , naturligtvis , europeiska standarder för livsmedelskvalitet inte tillämpas . - ( PT ) Jag förstår ledamotens oro fullkomligt och jag inser att det finns ett behov av vissa ansträngningar och en viss samstämmighet i frågan även inom Europeiska unionen .
Det är också viktigt att tänka på konsekvenserna framför allt vad gäller finansiering och ersättningar till jordbrukarna .
Denna fråga är dock , som ni känner till , i händerna på Europeiska kommissionen och kommer att utvecklas av kommissionen .
Rådets möjlighet att ingripa på detta område är begränsat . , rådet .
( PT ) Ärade ledamöter !
Dessa frågor går på djupet av den oro som ligger bakom det portugisiska ordförandeskapets program och den regering som tagit fram det .
Europeiska unionens råd är medvetet om problemen med de hemlösa och orsakerna är som ni vet många , från drogmissbruk till våld mot kvinnor och barn och långtidsarbetslöshet .
Det är ett extremt uttryck för sociala utslagning och fattigdom , som rådet försöker bekämpa på olika sätt .
Eftersom orsakerna är många måste förstås de olika politiska åtgärderna vara många och de måste diskuteras utifrån alla områden där unionen verkar och i hela den politik som kommer att bedrivas i denna fråga .
Det första politikområdet är kampen mot mäns våld mot kvinnor och barn , som många gånger leder till att kvinnorna flyr , med eller utan sina barn , och detta får ibland allvarliga konsekvenser för denna fråga .
Det kan också vara mäns och / eller kvinnors våld mot barn , vilket får barnen att fly , och som i dag leder till fenomen som drogberoende , prostitution etc .
För att bekämpa detta våld antog parlamentet och rådet i december Daphne-programmet , ett program för att bekämpa våldet mot kvinnor och barn och som snart kommer att inledas .
Detta program skall stödja de åtgärder som genomförs av icke-statliga organisationer inom detta område .
I början av maj i år kommer det portugisiska ordförandeskapet att anordna en konferens om våld mot kvinnor .
När det käller kampen mot narkotikamissbruk , är det lämpligt att erinra om programmet för förebyggande mot narkotikamissbruk antaget i december 1996 av Europaparlamentet och rådet i syfte att stimulera till ett arbete över olika politikområden och som framför allt beaktar de sociala och personliga konsekvenserna av detta problem .
Beträffande kampen mot arbetslöshet och social utslagning skulle jag vilja uppmärksamma , och detta har redan nämnts flera gånger här , dels av rådets ordförandeskap , dels av olika ledamöter , det initiativ Portugal har tagit till att i slutet av mars i år hålla ett extra europeiskt råd som ägnar sig just åt sysselsättningsfrågan , ekonomiska reformer och social sammanhållning , allt detta knutet till ett perspektiv av innovation och kunskap .
Det handlar om ett initiativ för att , som en av dess aspekter , bekämpa just den sociala utslagningen och för en social integrering genom att främja aktiva konkreta åtgärder och bättre samordning , dels av sysselsättningspolitiken , dels av en politik som kan bidra till en ökad europeisk konkurrenskraft och således öka utvecklingen av vår egen ekonomi med uppenbara effekter för förmågan att motverka alla de negativa sidoeffekter som den sociala utslagningen leder till och som givetvis är förbundet med fattigdom .
Vad gäller konkreta åtgärder för att bekämpa den sociala utslagningen vill vi påminna om att Europeiska kommissionen har meddelat att den kommer att lägga fram ett femårigt åtgärdsprogram i enlighet med artikel 137 i fördraget i syfte att bekämpa den sociala utslagningen .
Det portugisiska ordförandeskapet har redan tagit på sig att inleda arbetet så fort vi får kommissionens förslag .
Denna fråga , ärade ledamöter , och jag minns det på grund av mitt eget deltagande under senaste regeringskonferensen , aktiverade vissa europeiska länder under konferensen och som vi lyckades , kan vi säga , få in inom ramen för själva det reviderade Amsterdamfördraget .
Jag menar att detta ämne hela tiden måste finnas med , då det är en nyckelfråga där vi kan visa medborgarna den nytta de kan ha av Europa , i annat fall kommer det att bli svårt att uppamma någon vilja för mer Europa .
Men detta är ett problem , herr ledamot , som sträcker sig längre än det portugisiska ordförandeskapets sex månader .
Vi skall göra vad vi kan under dessa sex månader .
Herr talman !
Låt mig också välkomna rådets ordförande till kammaren .
Men jag tror inte att han svarade på min fråga som specifikt handlade om hur vi skall ta itu med hemlöshet och bostäder , och om det portugisiska ordförandeskapet kan tänka sig att på ett aktivt sätt föra ett samtal med de icke-statliga organisationer som är verksamma inom detta område .
Jag uppskattar och stöder fullständigt hans uttalande om behovet av flera strategier och ett sektorsövergripande förhållningssätt och också behovet av att bekämpa de underliggande orsakerna till utslagning , som kan leda till hemlöshet och omfatta drogberoende .
Min specifika fråga handlar om problemen med hemlöshet och om det nya ordförandeskapet kan ta nya initiativ för att försöka komma till rätta med en del av de svårigheter som rådsordföranden åsyftade vad gäller stöd på mellanstatlig nivå .
Jag anser att detta är ett område inom vilket Europa kan spela en mycket aktiv roll , även om det bara handlar om hur utbytet av erfarenheter och bästa metoder skall gå till mellan medlemsstaterna . - ( PT ) Herr ledamot !
När det gäller ordförandeskapets möjligheter att stödja de icke-statliga organisationernas arbete , särskilt när det gäller kampen för att lösa de personliga problemen för de hemlösa , vill jag säga att denna typ av initiativ är välkomna , och vi för vår del är öppna för att diskutera möjligheter att stödja dem .
Vi har samarbetat med de icke-statliga organisationerna i Portugal och angående några initiativ som dessa organisationer har presenterat inom ramen för det portugisiska ordförandeskapets verksamhet och som vi knyter till alla de angelägenheter som finns i vårt eget program .
Vi har inget specifikt konkret initiativ i denna fråga , vi är däremot inte låsta för tanken på att initiativ från de icke-statliga organisationerna som läggs fram för oss på detta område kan beaktas under vårt ordförandeskap .
Detta , vilket måste påpekas , inom ramen för det som hör till rådets verksamhetsområde .
Men vi måste förstå att allt det som handlar om kommissionens initiativrätt naturligtvis måste genomföras via kommissionen .
Herr rådsordförande !
Ni sade oss många saker om framtiden : vad kommissionen kommer att göra , vad ordförandeskapet kommer att göra i Lissabon m.m.
Och ni sade oss en sak som skrämmer mig , herr rådsordförande .
Ni sade att ni i Lissabon kommer att diskutera en utveckling som är mer dynamisk och konkurrensinriktad .
Jag blir rädd , herr rådsordförande , för det är en sådan utveckling som leder , åtminstone delvis , till social utslagning .
Jag kan inte förstå hur ni , med sådana åsikter , skall kunna ge ett svar på dessa problem .
Det som jag frågade och som jag frågar igen är följande : Vad är det portugisiska ordförandeskapets åsikt om de krav som kommer från t.ex. nätverken som bekämpar fattigdom och social utslagning , om fördelning av arbetstillfällen och social trygghet , om genomförandet av skattepolitiken , och då särskilt med avseende på det spekulativa kapitalet , om politiken för inkomstfördelning ?
Jag skulle vilja ha ett svar på frågan om det portugisiska ordförandeskapet har för avsikt att göra någonting vad beträffar dessa saker . - ( PT ) Herr ledamoten måste förstå att ett ordförandeskaps faktiska förmåga att vända på allmänna sociala eller ekonomiska tendenser under sin period är ganska begränsad .
Jag tycker att står helt klart att vår förmåga också är nära sammanbunden med vårt arbetsmetod med kommissionens initiativrätt .
Jag talade det extra Europeiska rådet och Portugals initiativ , jag talade också om framtiden för det finns ytterligare två sätt att se på frågan om social utslagning : ett av dem är de omedelbara åtgärderna som måste vidtas för att möta dess konkreta effekter , det andra är skapandet av förutsättningar för konkurrenskraft på ett internationellt plan så att vi kan förbättra det ekonomiska taket inom Europeiska unionen och få positiva sidoeffekter för problemen med social utslagning .
Det portugisiska ordförandeskapet har således inga universalmedel för att under sex månader lösa de frågor som vi alltid har med oss .
Vi är beredda att agera utifrån kommissionens förslag inom de områden som hör till gemenskapsbefogenheterna .
Vi har givetvis både möjlighet och intresse av att få i gång alla de åtgärder som läggs fram , framför allt av icke-statliga organisationer , men också i en traditionell mellanstatlig förbindelse på detta område .
Men vi måste vara medvetna om , herr ledamot , att det inte är möjligt att agera på ett område av så stor betydelse , ur ekonomiskt perspektiv , bara genom åtgärder som föreslås av ett ordförandeskap under en sexmånadersperiod .
Vi tycker därför att det är klart att alla de åtgärder vi har pekat på angående strategier på längre sikt , oberoende av att vi vet att en del av de hemlösa på lång sikt kan vara döda , är de som kommer att göra det möjligt att få en hållbar politik i Europeiska unionen .
Det är dessa strategier som vi vill försöka bidra till på bästa möjliga sätt under vårt arbete .
Fråga nr 12 från ( H-0801 / 99 ) Angående : Portugals ordförandeskap och utvecklingspolitiken Kommer rådets sittande ordförande att uttala sig om prioriteringarna för Portugals ordförandeskap när det gäller utvecklingspolitiken , Lomékonventionen och hanterandet av svältsituationer ? , rådet .
( PT ) Herr talman !
Frågan om den europeiska politiken för utvecklingsbistånd är en fråga som har genomgått en påtaglig utveckling de senaste åren .
Vi deltar särskilt i all debatt om förnyandet av Lomékonventionen och fastställandet av den nya avtalsram som skall efterträda Lomékonventionen .
Jag anser att detta är några frågor - och jag säger det med myndigheten hos den som har deltagit i förhandlingarna , dels när Portugal gick med i Lomé III , dels som ordförande för den portugisiska delegationen i förhandlingarna om Lomé IV - som allmänheten och särskilt regeringarna ( och även ledamöterna här ) genomgående vill ha svar på , det vill säga hur effektiva de anslag som har getts i utvecklingsbistånd har varit i kampen mot de negativa aspekter de har varit avsedda för .
Det portugisiska ordförandeskapets prioritering kommer att vara att under januari månad genomföra ett informellt möte med utvecklingsministrarna vilket skall ligga till grund just för att fastställa en europeisk strategi för utvecklingssamarbetet .
Vi anser alltså att det är mycket viktigt att framför allt inom OECD : s kommitté för utvecklingsbistånd och i den allmänna ramen för förberedelser för nästa UNCTAD , kunna ha en kollektiv ståndpunkt och organiserad så att vi får en idé om hur unionens resurser för utvecklingsbistånd används .
Varför det ?
Detta också därför att våra egna nationella parlament är uppmärksamma , precis på samma sätt som detta parlament måste vara på ett gemenskapsplan , hur dessa anslag tilldelas och används .
Vi är angelägna om att se till att denna diskussion kan vara användbar , fruktbar och få konkreta resultat , framför allt i vår framtida verksamhet på ett internationellt plan .
Vi tycker också att vår nya avtalsmodell som definieras av Lomékonventionen är en mer ansvarsfull , balanserad och effektiv modell än i de tidigare Yaoundé- och Lomékonventionerna .
Jag skulle också vilja säga , herr talman , ärade ledamöter , att i hypotesen om att ännu kunna genomföra toppmötet mellan Europeiska unionen och de afrikanska länderna , är naturligtvis frågorna om utvecklingssamarbete , och en allmän tolkning av hur utvecklingsfrågorna kan behandlas inom ramen för bilaterala förbindelser mellan dessa två områden , centrala för vår inriktning och kommer att utgöra ett av de centrala ämnena för denna dagordning .
Jag vill tacka ordförandeskapet för det omfattande svaret på min fråga , och även ministern som uttalade sig i utskottet för utveckling och samarbete förra veckan i Bryssel , där han presenterade ståndpunkten .
Men det finns fortfarande vissa frågor som är obesvarade .
Det verkar inte finnas någon betoning på kampen mot aids i programmet. aids-situationen i Afrika är nu så allvarlig att det dör fler människor i aids än p.g.a. krig .
Jag hoppas att ministern kommer att lägga ned en viss tid på denna specifika fråga .
Det finns tillgängliga mediciner i Förenta staterna , men Förenta staterna tillverkar dem inte tillräckligt billigt för de drabbade i Afrika .
Jag vill fråga ministern vad han tänkt göra åt situationen som håller på att utveckla sig i Etiopien , där det råder torka , där skörden har slagit fel och där vi om sex månader oundvikligen kommer att vara tillbaka i det läge som rådde för några år sedan i landet , med svält och tusentals människor som dog .
Samtidigt är det krig mellan Eritrea och Etiopien och vapenindustrin i Europa är inte sen att skicka vapen , efter vilka vi skickar bröd . - ( PT ) Ledamoten måste förstå att jag först och främst inte håller med om er tolkning av min kollegas inlägg under mötet med utskottet för utveckling och samarbete , det finns inget motsägelsefullt mellan dessa ståndpunkter , snarare tvärtom .
Vi kan inte i ett ordförandeskapsprogram , så vitt vi inte drabbas av storhetsvansinne , göra ett uttömmande inventarium av all möjliga och imaginära situationer för alla stora frågor som dyker upp inom ramen för internationella förbindelser .
Det skulle som ni förstår vara enkelt att göra det .
Det räcker med att ta en ordlista över utveckling och placera dem där , ord efter ord .
Vi är tillräckligt ansvarsfulla att förstå att vi bara kan ta upp de vi har förutsättningar att klara av under vårt ordförandeskap och inom vilket - och vi bör alltid vara medvetna om detta - regeringarnas kapacitet inom rådet .
Vi bör inse att det finns begränsningar vad gäller förvaltningen av de nationella vägledande programmen .
Ledamoten tog upp frågan om Etiopien , vilken hör till de nationella orienteringsprogrammen , men det finns som ni känner till olika gemenskapsåtgärder till kampen mot Aids , och i denna aspekt har ni rätt , herr ledamot , troligen agerar inte heller USA på bättre sätt .
När det gäller politiken för utvecklingsbistånd anser jag att Europa inte har något att oroa sig över av det enkla skälet att vårt agerande i denna fråga kan mäta sig med USA : s .
Ledamotens fråga kom in på frågan om rustningsproblemets effekter , och det är en mer långtgående politisk fråga som jag inte tycker inryms i denna fråga men som rådet naturligtvis i framtiden kommer att ta itu med , om man anser att man skall det , och lösa genom att sätta in det i sitt speciella sammanhang .
Är rådet medvetet om de sociala problem som den EU : s livsmedelsexport till u-länderna som sker till priser under produktionskostnaderna ?
Har ordförandestaten för avsikt att göra någonting åt den saken ? - ( PT ) Fru ledamoten tar upp ett traditionellt problem inom livsmedelsbiståndet , det vill säga , om livsmedelsbiståndet leder till nedgång för jordbrukarna i utvecklingsländerna .
Detta är en återkommande fråga som aldrig har fått något svar inom området för utvecklingsbistånd och som traditionellt ställs eftersom många åtgärder beträffande livsmedelsbistånd i själva verket har negativa effekter för förmågan att skapa jordbruksstrukturer i dessa länder och främst för familjejordbruk .
Jag har inte lösningar på detta och efter mina dryga tjugo års erfarenheter av dessa frågor tror jag inte att har det .
Eftersom frågeställaren är frånvarande , bortfaller fråga nr 13 .
Frågorna nr 14 , 15 och 16 kommer på begäran av rådet att tas upp tillsammans , trots att de behandlar skilda ämnen : Fråga nr 14 från ( H-0809 / 99 ) : Angående : Europeisk kultur Begreppet Europa har en i grunden kulturell innebörd .
Och Europeiska unionen kommer att etablera sin ställning och väcka gensvar över världen om den visar att en av dess grundläggande prioriteringar är den kulturella dimensionen , i förening med den ekonomiska .
Det är beklagligt att man inte är tillräckligt medveten om det faktum att även kulturen är en stor ekonomisk tillgång .
Därför får kulturen också bara futtiga anslagssummor och även de verkar vara på väg att försvinna för rådets och kommissionens del .
Detsamma gäller tyvärr även för den andra stora ekonomiska tillgången - idrotten .
Om man utnyttjade idrotten på ett lämpligt sätt skulle den kunna bli till stor hjälp för att ta itu med EU : s huvudproblem , dvs. arbetslösheten , och även se till att det flödar in extrainkomster från det internationella utnyttjandet .
På det sättet har USA dominerat världsmarknaden för musik och underhållning , och genom detta framför allt yngre generationers tänkande , preferenser och bildning .
Är rådet berett att vid regeringskonferensen medge att även kulturen är en ekonomisk tillgång och prioritera den på motsvarande sätt ?
Fråga nr 15 från ( H-0814 / 99 ) : Angående : Europeisk sysselsättningspolitik Har rådet för avsikt att inför regeringskonferensen utforma en europeisk sysselsättningspolitik som är försedd med tillräckliga budgetmedel och som tar hänsyn till att det enligt unionens officiella statistik finns ett direkt samband mellan arbetslöshet och låg produktivitet ?
Fråga nr 16 från ( H-0005 / 00 ) : Angående : Rådets ordförandeskap Ordförandeskapet i EU roterar för närvarande mellan medlemsstaterna enligt ett system som Europeiska rådet enats om .
Med tanke på att en ny regeringskonferens snart inleds verkar det nu lämpligt att se över systemet .
Förenade kungarikets konservativa ledamöter i Europaparlamentet anser att den medlemsstat som innehar ordförandeskapet skall utgöra ett ytterst gott exempel ifråga om införlivandet av EU : s lagstiftning till nationella lagar och efterlevnaden av EU : s lagstiftning då den trätt i kraft .
Kan rådet med anledning av detta vid regeringskonferensen diskutera ett annat system med vilket man garanterar att en medlemsstat endast kan bli ordförandeland om det uttryckligen visar tillräcklig respekt för EU : s lagar ?
Kan rådet dessutom kommentera förslaget att den medlemsstat som ligger i nedre delen av en " topplista " över införlivandet av direktiv och antal fall anmälda till EG-domstolen , skall avstängas från ordförandeskapet i Europeiska unionens råd ? , rådet .
( PT ) Låt mig beträffande Marinos frågan , för det första understryka det faktum att rådet är helt medvetet om att den kulturella dimensionen utan tvivel är en av de främsta triumferna för Europa och att vi måste uppbåda alla våra krafter för att skydda vår kulturella identitet .
De här sakerna har funnits med på flera olika sätt i unionens bekräftelse utåt och främst inom ramen för de angelägenheter vi har haft inom Världshandelsorganisationen .
Rådet underskatter inte heller betydelsen av kulturen och idrotten på ett ekonomiskt plan .
Tillåt mig därefter , herr ledamot , att uppmärksamma det faktum att , om den kulturella dimensionen i den europeiska politiken bör uppmärksammas av behöriga myndigheter , bör detta i princip ske under subsidiaritetsprincipens beskydd , med tanke på det som bör genomföras på såväl nationell nivå som på gemenskapsnivå .
När det gäller Nogueira Románs fråga , om sysselsättning , hänvisar jag till vad jag sade nyligen : denna fråga är fortfarande en fråga som oroar medlemsstaternas ledamöter och regeringar och kommer givetvis att vara en central angelägenhet för det portugisiska ordförandeskapet .
Det finns till och med de som säger att den är för central för det portugisiska ordförandeskapet , med tanke på att Portugal inte ens till de länder som har en hög arbetslöshet , men vi har ett europeiskt perspektiv på hur vi skall utöva vårt ordförandeskap .
Jag tror att Europeiska rådet i Lissabon och genomförandet av det jag nämnt tidigare svarar perfekt mot detta .
Jag anser , herr talman , att de frågor ni har ställt hör ihop med frågorna från ledamöterna Bushill-Matthews och Nogueira Román .
Jag skulle vilja säga angående den kommande regeringskonferensen att rådet bara kan hänvisa ledamöterna till slutsatserna från Europeiska rådet i Köln och i Helsingfors , vilka fastställde mandaten för denna konferens , och följa åliggandena för själva konferensen , som har en mellanstatlig struktur , och inom ramen för sitt mandat , analysera i vilken mån de frågor som ställts av ledamöterna kan behandlas under konferensen .
Men naturligtvis kommer den breda tolkning det portugisiska ordförandeskapet ämnar göra av Europaparlamentets ledamöters roll i den förberedande gruppen att tillåta dem att komma med inlägg och kanalisera det som parlamentet är angeläget om i den förberedande gruppen .
Givetvis kommer också Europaparlamentets talman att ha möjlighet att på ministernivå lägga fram dessa frågor .
När det gäller de halvårsvisa ordförandeskapen handlar det om en fråga som inte det portugisiska ordförandeskapet tänker ta upp som initiativ under den kommande regeringskonferensen .
Om någon vill ta upp det noterar vi det och underställer det konferensen .
Jag tackar rådsordföranden och framför till honom min personliga välkomsthälsning till den portugisiska regeringens ordförandeskap .
Tillåt mig att tala om för honom hur vältalig och kunnig han är om de europeiska frågorna .
Dock gav han tyvärr inte i mitt eget ärende ett svar som jag skulle kunna finna tillfredsställande .
Eftersom rådet erkänner kulturens stora betydelse som ekonomisk handelsvara , borde det , enligt min åsikt , visa det även i praktiken .
Och jag är rädd för att ursäkten att kultursektorn styrs av subsidiaritetsprincipen , och följaktligen är de nationella regeringarnas ansvar , är ett svepskäl .
För den fråga som jag ställde och som förblev obesvarad är varför rådet , liksom för övrigt också kommissionen , när Europaparlamentet begär ökade anslag för att finansiera Europeiska unionens kulturprogram , regelmässigt minskar dessa och ibland till och med avslår dem helt .
Det visar i praktiken rådets ointresse för kulturen , trots rådets motsatta försäkringar om att det tillskriver kulturen stor betydelse .
Jag skulle alltså vilja fråga rådet om det är berett att från och med nu stödja kulturen , med samma iver som det subventionerar bananerna , humlen , korna och cannabisen . - ( PT ) Vi har inte , herr ledamot , ett ekonomistiskt koncept för vårt utövande av det portugisiska ordförandeskapet och därför ligger den kulturella dimensionen som ni förstår i centrum för vårt arbete .
Men dessa kulturella dimensioner har nästan alltid i sig en ekonomistisk egenskap , det vill säga , de medel som kan mobiliseras just för att stödja de kulturella åtgärderna .
Detta är en dimension det är svårt att komma förbi inom Europeiska unionens område och framför allt inom ramen för rådet .
För vår del kommer vi att försöka stärka och befästa den europeiska ställningen vad gäller kulturell egendom och verksamheten inom detta område eftersom vi anser att detta är en viktig identitet för unionens egen bild och unionens specifika identitet .
Det är och kommer i framtiden att vara knutet till vad som sker inom ramen för Världshandelsorganisationen .
Denna fråga har som ni vet för vår del och för rådets del behandlats på lämpligt sätt och det var framför allt möjligt att finna ett uttryck i linje med det mandat kommissionen fått för förhandlingarna inom nästa runda i Världshandelsorganisationen , där denna fråga är central .
Jag skulle dock vilja tillägga att när det gäller kulturpolitiken , och främst det audiovisuella området , kommer det portugisiska ordförandeskapet att verka för en särskild uppmärksamhet på att fördjupa och berika den europeiska audiovisuella politiken genom antagandet av ett Media-Plus-program som skall kunna motsvara de stora europeiska intressena .
Vi avser också att inleda en ny mer innovativ debatt , i frågan om det europeiska kinematografiska arvet , då vi anser att detta måste vara en av de viktigaste beståndsdelarna i en europeisk kulturell identitet och en europeisk audiovisuell ekonomi .
Ordförandeskapet kommer även att koncentrera sig på diskussionerna om att införa ett system för digital-TV i Europa , vilket kommer att vara föremål för en konferens som vi kommer att arrangera under det portugisiska ordförandeskapet , tillsammans med kommissionen , i februari 2000 .
Men kulturen , herr ledamot , i Europeiska unionen är en fråga som ständigt dyker upp på regeringskonferensernas dagordningar .
Om bara det som definieras som den femte förhandlingsdelen under den kommande regeringskonferensen kunde uppnå enighet om att inkludera det kulturella området , skulle detta kunna föreslås , dels av medlemsstaterna , dels av Europaparlamentets ledamöter som kommer att delta i den förberedande gruppen .
Naturligt skulle det kunna vara ett framsteg om denna fråga kunde uppnå enighet inom ramen för regeringskonferensen .
Det återstår att se om det finns en enighet om detta eller ej .
Därefter får vi ser .
För vår del kommer vi att ta notis om de förslag som lagts fram i detta ämne .
Herr talman !
Låt mig instämma i övriga talares önskan om att Portugal skall få ett framgångsrikt ordförandeskap .
Jag lade märke till att ni sade att denna specifika fråga för tillfället inte fanns på er dagordning för nästa regeringskonferens , men om man önskade detta skulle ni överväga att ta med den .
Nu är det så att jag och mina 35 brittiska konservativa kolleger önskar detta och vill att ni skall överväga det .
Jag har förståelse för att det är en utmanande fråga .
Den är avsedd att vara utmanande , eftersom detta är en mycket allvarlig fråga då vissa länder inte respekterar EG-lagstiftningen i tillräcklig omfattning .
Vi måste hitta ett sätt utöva påtryckningar på dessa länder så att de gör det , så att vi och medborgarna återigen kan känna en gemenskap .
Jag kan inte komma på ett bättre sätt att göra det .
Kan ni ? - ( PT ) Frågan är om den europeiska dimensionen kommer att förstärkas mer eller mindre genom att den integreras i fördragen .
Detta är en fråga som måste behandlas på regeringskonferensen , som ni förstår , och det är ett av de ämnen som bara ett extra europeiskt råd kan bevilja det portugisiska ordförandeskapet att följa upp , eftersom frågan ligger utanför den institutionella ram inom vilken den kommande regeringskonferensen kommer att genomföras .
Nu är regeringskonferenserna en slags händelse och det kan också bli en slags julgran .
Därför kan man inte utesluta möjligheten att dessa återkommande frågor , och som har passerat konferens efter konferens , kan tas upp .
Problemet är om vi kan uppnå enhällighet i detta ögonblick , inom ramen för Europeiska unionen , för att denna fråga skall tas upp , särskilt med tanke på att om denna typ av fråga tas upp , kommer troligen andra liknande frågor att utöka konferensens dagordning .
Ordet går till Dimitrakopoulos för en ordningsfråga .
Jag ber er att fatta er kort . )
Herr talman !
Jag förstår att jag måste fatta mig kort .
Jag tyckte mycket om det som Seixas da Costa sade om jultomten .
I Spanien skickar vi brev till de tre vise männen .
Jag vill bara påminna er om att Europaparlamentet redan har skickat sitt brev med betänkanden till de tre vise männen .
Nu är det ordförandeskapet och rådet som måste komma med de presenter vi bett om i brevet .
Som jag misstänkte så var det inte en ordningsfråga det var frågan om , utan en avrundning på debatten .
Vi tackar Seixas da Costa , men han kan också skriva ett brev till de tre vise männen . - ( PT ) Jag vill bara säga att denna fråga av julkaraktär som ledamoten har tagit upp är av största vikt .
Bara det att i detta fall har jultomten någon som bestämmer och således kan jultomten bara ge presenter när han ges tillstånd av andra att göra det .
Det hänger inte på det portugisiska ordförandeskapet att ge de presenter som alla vill ha , och speciellt de som Europaparlamentet vill ha .
Efter denna intressanta åsiktsyttring , och i enlighet med arbetsordningen , besvaras frågorna nr 17 till 27 skriftligen .
Jag förklarar härmed frågestunden till rådet avslutad .
 
Kapitalskatt Nästa punkt på föredragningslistan är gemensam diskussion om följande punkter : den muntliga frågan ( B5-0004 / 2000 ) från Désir m.fl. till rådet om rådets synpunkt på idén om en kapitalskatt den muntliga frågan ( B5-0005 / 2000 ) från Désir m.fl. till kommissionen om kommissionens synpunkt på idén om en kapitalskatt .
Fru talman , herr rådsordförande , herr kommissionär !
Alla kunde i samband med Asienkrisen 1997 , eller krisen i Mexiko 1995 , eller det europeiska monetära systemet 1993 , notera de skador som ekonomisk spekulation kan leda till på ekonomin i ett helt land , särskilt när denna utövas mot valutorna .
1 500 till 2 000 miljarder euro växlades varje dag på finansmarknaden , vilket på tre eller fyra dagar motsvarar världens hela årsproduktion , världens BNI , om ca 6 000 miljarder euro .
Detta innebär att största delen av dessa finanstransaktioner är rent spekulativa , utan koppling till handel med varor eller till investeringar .
Men en felaktig förflyttning av dessa avsevärda belopp kan på några timmar leda till att en valuta eller ett lands ekonomi rasar samman , och tvinga hela landets befolkning ned i en tillbakagång .
Inför denna situation har man visat nytt intresse för förslaget från nobelpristagaren James Tobin om att inrätta en skatt på transaktioner med valutor , som skulle vara mycket låg , så att den inte skadar handeln med varor eller investeringarna , men fungerar som ett gruskorn i spekulationens maskineri , dvs. bromsar det ökande antalet kortsiktiga transaktioner .
Märk väl att detta förslag till skatt , som förefaller orsaka så starka känslor hos vissa , skulle vara världens lägsta skatt , den lägsta i världens skattehistoria , men den skulle också vara ett sätt att återerövra de demokratiska områden som finansvärlden lagt beslag på .
En anledning till att förslaget rönt framgång , liksom kampanjerna från de icke-statliga organisationerna såsom ATTAC , Solidar eller andra som populariserat det , är också att det skulle lösgöra resurser för utvecklingsprogram i de fattigaste länderna , inom utbildnings- eller hälsoområdet .
Det är en slags omfördelning i en värld där det både finns allt fler rika och allt fler fattiga .
Ett stort antal personer och institutioner har yttrat sig positivt för denna skatt , såsom Brasiliens president , Fernando Cardoso , Finlands regering , Canadas parlament i mars förra året , men också Lionel Jospin redan 1995 .
Förslaget har diskuterats i flera nationella parlament i Europeiska unionen .
Svaret har ofta varit att frågan inte endast kan behandlas på nationell nivå och Europeiska unionen är rätt forum att ta upp frågan i , vilket är anledningen till den muntliga frågan till rådet och kommissionen som vi lämnat in tillsammans med 37 andra parlamentsledamöter .
Jag gläds åt förslaget till kompromissresolution , som vi uppnått tillsammans med GUE-gruppen , Gruppen De gröna , den liberala gruppen och PSE-gruppen , och där vi ber kommissionen att lägga fram en rapport till parlamentet inom sex månader om genomförbarheten av denna skatt samt granska de ekonomiska påtryckningar och sanktioner som skulle kunna tillämpas mot de länder som uppmuntrar skatteflykt eller underhåller skatteparadis .
Man invänder ofta att en sådan skatt skulle kringgås , men det kan man säga om alla skatter och om man hade lyssnat på det argumentet skulle vi aldrig ha infört någon skatt .
I resolutionsförslaget krävs också att man före nästa årsmöte i Internationella valutafonden lägger fram ett dokument om den ståndpunkt som utarbetats av kommissionen och rådet .
Jag tror att Europeiska unionen måste ta initiativet , att den också , såsom krävs i förslaget till resolution , skall föreslå detta initiativ till G7-länderna eftersom det i första hand är en politisk fråga .
Om unionen tar initiativet drar det andra med sig , eftersom debatten äger rum överallt , inbegripet Förenta staterna och Japan , och det finns en allt starkare strävan i världen efter att den skall styras inte av handlare utan av medborgare , deras parlament , regeringar och demokratiska institutioner .
Jag tror att Europa måste spela en roll i denna nya internationella reglering och jag är mycket glad över att frågan , genom denna debatt och förslaget till resolution , finns på dagordningen för den europeiska integrationen . , rådet .
( PT ) Fru talman !
Jag har inte mycket att komma med i denna fråga .
Rådet har hittills inte diskuterat möjligheten att införa en skatt på kapitalrörelser , så som professor Tobin har föreslagit .
Det handlar om ett kreativt initiativ , som vi vet har tagits emot väl inom diverse sektorer på internationell nivå och i olika politiska sektorer i Europa , men det är en fråga som det inte har kommit några förslag eller initiativ om från kommissionen .
Då det tillkommer kommissionen att ta eventuella initiativ kan inte rådet ta ställning i denna fråga . .
( NL ) Fru talman !
Inkomstgrunden för Tobinskatten skulle bestå av mycket korta valutatransaktioner .
Sådana transaktioner , heter det , har mycket litet samband med grundläggande ekonomiska variabler .
Det betonade också Désir alldeles nyss .
Förespråkarna , som till exempel Désir , menar då också att en internationellt tillämpad Tobinskatt i princip skulle minska de spekulativa transaktionerna och alltså även valutakursernas nyckfullhet och det skulle leda till en förbättrad ekonomisk välfärd .
Med tanke på den stora omfattningen av de korta ekonomiska flödena skulle till och med en Tobinskatt med lågt nominellt värde ge rejäla skatteinkomster .
I verkligheten var skälet till det ökade intresset för Tobinskatten och för andra internationella finanskällor i mitten på nittiotalet inte av ekonomisk art .
Det var nämligen den skattens möjlighet att skapa inkomster för offentliga internationella program i en tid då efterfrågan på sådana fonder ökade snabbt och det blev allt svårare att finansiera dem .
Nyligen konstaterade kommissionen ett pånyttfött intresse för en global skatt som till exempel Tobinskatten som medel för att uppnå en , skulle man kunna säga , socialt försvarbar globalisering .
Även Désir har nämnt det växande intresset från olika håll .
Om Tobinskatten ensidigt skulle tillämpas för att hindra angrepp mot en viss valuta så skulle den här skatten inte kunna vara effektiv och den skulle då kunna skada den finansiella inhemska marknaden .
Ännu värre , på lång sikt är det möjligt att Tobinskatten undviks för flera fonder genom att utländska valutatransaktioner överförs till finansiella centrum off-shore .
I det fallet skulle skatten kunna leda till en nettoförlust i totalekonomisk välfärd .
Tobinskatten kan alltså endast fungera om tillräckligt många industriländer är villiga att delta .
Även om Tobinskatten utformats för att stävja valutaspekulationerna så finns fortfarande risken att även andra flöden än de spekulativa drabbas och det är inte meningen .
Av dessa skäl ser jag ingen anledning till att införa en europeisk Tobinskatt .
Kommissionen är i alla fall motståndare till varje försök att begränsa kapitalrörligheten i Europeiska unionen .
I den mån den åtgärden skulle kunna ses som en indirekt begränsning av kapitalflödet skulle den strida mot Romfördraget .
Rätt sätt att handskas med spekulationer , tycker jag , är att avlägsna de verkliga orsakerna till finansiell förvirring och inte att försöka undertrycka symptomen genom att införa hinder för marknadernas funktion .
Fru talman , herr kommissionär , mina damer och herrar !
Jag måste ännu en gång säga några saker med anledning av det förfaringssätt och den ideologiska taktik som lett fram till den här muntliga utfrågningen .
Jag gör det också eftersom jag vet att vår kritik delas av många socialdemokrater i kammaren , och inte bara av de ekonomisk- och finanspolitiska experterna .
Vi känner till problemet .
Det är marknadernas instabilitet till följd av spekulationer .
Men förslagsställarna måste få veta att det inte är varje instabilitet som är en följd av spekulationer - vilket också kommissionären med kraft redogjort för .
Tobinskatten skulle varken ha kunnat förhindra kriserna i Europeiska ekonomiska samarbetsområdet ( EES ) år 1992 och 1993 eller kriserna i de sydostasiatiska valutorna år 1997 .
Initiativtagarna till denna utfrågning föreslår ingen lösning utan ropar efter nya föreskrifter , mer byråkrati , efter åtgärder mot marknadsmekanismerna och tillskriver plenumet en intergroup-uppfattning ; samtidigt utestänger de det ständiga parlamentariska utskottet vilket står i motsättning till flera parlamentsbeslut .
Utfrågningen är som jag ser det tydligt ideologiskt motiverad och inte inriktad på att nå en lösning .
Jag anser att detta är fel väg av flera anledningar .
Vad är anledningen till att vi motsätter oss Tobinskatten och anser den vara så betänklig ?
För det första för att den skulle innebära en stark belastning på kapitalmarknaderna , vilket även kommissionären bekräftat .
Även en mycket blygsam skatt skulle få allvarliga följdverkningar på kapitalmarknaderna , eftersom en sådan spekulationsskatt i hög grad skulle reducera räntabiliteten på investeringarna .
Dessutom skulle en sådan åtgärd också få en stark påverkan på finansmarknadernas utveckling .
Det skulle stå i motsättning till principen om fria kapitalrörelser , som är en central del i den inre marknaden .
För det andra : Spekulationskapitalet är svårt att identifiera .
För det tredje : Skattemässiga åtgärder kan lätt kringgås om de inte införs i alla länder - i annat fall blir det för många kryphål .
För det fjärde : Åtgärden är tekniskt sett så gott som ogenomförbar ; den skulle leda till mycket byråkrati , förvaltning och okontrollerbara skeenden .
Den åtgärd vi bör vidta ingår som en del i resolutionen som vi har här i dag .
Det handlar om stärkt bankkontroll .
Det handlar om klargörande av var ansvaret för transaktioner ligger .
Det handlar om ramar för reglering på internationell nivå .
Det handlar om kontroll av nationella gränser med avseende på om de stämmer överens med Baselkommitténs regler och hur dessa kan spridas i ökad mån .
I föreliggande resolution har jag hittat ett stort problem på en central punkt , ett problem som vi inte kan acceptera i dess nuvarande form .
Det gäller punkt 9 .
När vi nu har lyssnat på vad kommissionären har sagt vet vi att kommissionens sakkunskap kommer att leda till ett nej till Tobinskatten .
Om nu sakkunskapen , debatten och argumenten ligger i linje med vår beskrivning - vilket jag tycker - så är det oansvarigt av kommissionen att utfärda en bestämmelse för ytterligare sex månader vilket medför osäkrare förhållanden på finans- och kapitalmarknaden .
Kapitalmarknaden behöver inte osäkrare förhållanden från vår sida , utan tydlighet .
Vi avvisar därför punkt 9 och kräver delad omröstning .
Fru talman !
Debatten om beskattning av kortfristiga finansiella transaktioner är inte ny .
I tjugo år har vi diskuterat förslaget om Tobinskatt ; men trots det är frågan alltid aktuell och vi behöver verkligen konkreta och redliga svar på grundfrågan utifrån noggranna studier .
Vi måste få reda på hur önskvärt och görligt det är att beskatta de kortsiktiga finansiella transaktionerna .
Frågan infinner sig i dag också faktiskt i en annan dimension , med tanke på att 1 500 miljarder US-dollar dagligen dygnet runt jagar efter attraktiva investeringar , varav högst 3 procent har samband med den reella ekonomin .
Vi engagerar oss visst i finansmarknadernas stabilitet - inte för finansmarknadernas skull utan för vår egen , eftersom det handlar om vår tillväxt , våra investeringar och våra arbetstillfällen i Europeiska unionen .
Här måste vi fråga oss vilka instrument vi kan använda för att skapa en viss ordning som hittills faktiskt saknats .
Vi har själva medverkat till avregleringen av systemet med finansiella transaktioner , men vi har ännu i dag inget fungerande regelverk och det har vi bittert fått erfara i samband med efterverkningarna av kriserna i Asien och Latinamerika .
Därför är det hög tid att vi börjar tänka dels på kontrollregler och dels på öppenhet på finansmarknaderna och deras informationsflöde .
Det är viktigt att vi vet vilka aktörerna är och vilket rykte de har .
Vi måste också fråga oss om vi inte är förpliktade att verka för skattemässig rättvisa .
I en tid när skattebelastningen av arbetet som produktionsfaktor stiger i hela Europa - liksom även internationellt sett - måste vi överväga hur vi kan åstadkomma en effektiv beskattning av kapitalvinster ; då måste vi även ställa frågan om beskattning av kortsiktiga finansiella transaktioner .
Jag menar att det är helt nödvändigt att vi får en grundlig rapport med slutsatser från kommissionen ; då kan vi i Europaparlamentet undersöka om vi inte måste se till att Europeiska unionen tillsammans med USA och Japan bestämmer sig för att åstadkomma en internationell solidaritet i syfte att ekonomin och finansmarknaderna skall bli stabilare och säkrare .
Det är denna intention som står bakom den muntliga utfrågningen ; vi i parlamentet har sedan att inom ramen för betänkandena i de ordinarie förfarandena via utskotten och plenarsammanträdena åstadkomma ett balanserat och framtidsinriktat förslag . )
Fru talman , ärade kollegor !
Å Europeiska liberala , demokratiska och reformistiska partiets grupp vill jag säga att jag förvånas över den debatt som nu sysselsätter oss om internationella kapitalflöden och en eventuell beskattning som , även om det inte nämns i texten , verkar vara ett försök att återuppliva Tobins förslag om beskattning , som lades fram för några år sedan och som vår grupp kraftfullt motsatte sig under den föregående mandatperioden med en rad klara och tydliga argument presenterade av ordförande Cox .
Argument som jag blygsamt verkar vara tvungen att upprepa , eftersom samma fråga på nytt dyker upp .
Vi motsätter oss en sådan beskattning , om den nu kan genomföras , eftersom den inte skulle tjäna de syften som Tobin förespeglade och som vänstern i kammaren verkar vilja återuppliva .
För det första finns det inga bevis på att en beskattning av det internationella kapitalflödet skulle kunna minska instabiliteten på de internationella marknaderna .
Tvärtom , eftersom inte alla länder kommer att acceptera det , skulle vi bana väg för spekulation och bedrägeri vilket skulle förorsaka förgänglighet , instabilitet , osäkerhet , dunkelhet och illojal konkurrens för de finansiella tjänster som är verksamma på en internationell nivå .
Idén med att erhålla medel för länder som är i behov av ekonomiskt stöd är dessutom mycket komplicerat , när man nu tänker på hur det hela skall tillämpas i praktiken , vilket gör det fullständigt omöjligt .
Ärade kollegor , den här debatten är falsk och fyller inte något annat ändamål än att täcka en politisk målsättning , en målsättning utan grund och tekniskt ogenomförbar .
Dessutom - nu när vi befinner oss här i Europaparlamentet - om vi inte har lyckats träffa en överenskommelse om de skatteåtgärder som kommissionen föreslår för Europeiska unionen , hur har vi då tänkt nå en skatteöverenskommelse på internationell nivå .
Jag antar att de kommer att säga : Få se om ni först har förmåga att nå en skatteöverenskommelse inom unionen !
Ärade kollegor , Liberala gruppen har inte velat stänga dörrarna för en ny analys av frågan och därför har vi i det gemensamma resolutionsförslaget accepterat att en studie genomförs om möjligheten och fördelarna med nämnda beskattning av vissa delar av det internationella kapitalflödet .
Jag är säker på att studien - om den genomförs objektivt och med kännedom om den finansiella marknaden och dess mekanismer på internationell nivå - kommer att visa att det varken är lämpligt eller möjligt , inte bara när det gäller tillämpningen utan också som medel för att uppnå de mål som eftersträvas .
Globaliseringen är i sig positiv .
Aldrig någonsin har ekonomin vuxit så snabbt och globalt gynnat så många länder .
Anledningen är ett progressivt öppnande och en ökad frihet när det gäller utbyte av varor och tjänster på internationell nivå samt större kapacitet för att det skall finnas lämpliga kapitalflöden .
Analysera den ekonomiska utvecklingen under de senaste åren , och är ni objektiva så kan ni av resultatet själva konstatera att den inte styrts av någon politisk inriktning eller färg .
Som sagt så motsätter vi oss inte att studien genomförs .
Vi stöder övergångsresolutionen så att studien kan göras , men eftersom den också finns med i resolutionsförslaget vidhåller vi att det är just genom en avreglering och ett internationellt öppnande som vi kan få ekonomisk tillväxt , såväl på nationell som internationell nivå .
Fru talman , herr kommissionär !
Jag tror inte problemet är att ideologisera debatten utan att bedriva politik .
Jag tror att man , såsom Randzio-Plath sade , måste erinra om att anledningen till att ett antal parlamentariker önskar ta upp frågan igen är de senaste internationella finanskriserna och deras ekonomiska , sociala och miljömässiga konsekvenser i en rad länder , något som alla känner till .
Den huvudsakliga målsättningen med denna diskussion är att se vilka instrument den internationella gemenskapen kan förfoga över för att stabilisera det internationella valuta- och finanssystemet .
Herr Bolkestein !
Ur den synvinkeln isolerar förslaget till resolution inte frågan om Tobinskatten .
Om ni läser det noggrant är detta förslag till skatt på kapitalflödet ett instrument bland andra , för att försöka tvinga de internationella investerarna till ett ansvarsfullt uppträdande på finansmarknaderna .
För det andra sägs inte i resolutionen att vi vill ha ett initiativ på enbart europeisk bas .
Det är anledningen till att vi uttryckligen hänvisar till höstsammanträdet i Internationella valutafonden för att Europeiska unionen , dvs. kommissionen , men också rådet , skall inta en ståndpunkt om hur de kommer att försvara möjligheten att stabilisera det internationella finans- och valutasystemet , och införa en internationell beskattning .
Jag vill inte att det skall föreligga några missförstånd i debatten .
Vi miljöpartister vill inte ha en alibiresolution .
Det handlar inte om att lägga ytterligare en studie till det tiotal som redan genomförts - kommissionens skulle säkerligen vara intressant - utan om att från kommissionen och rådet , dvs. från varje regering som unionen består av , erhålla en tydlig , positiv eller negativ politisk ståndpunkt , om de är beredda att i berörda allmänna sammanhang dvs .
Internationella valutafonden till att börja med , försvara möjligheten med en sådan skatt jämfört med andra nödvändiga instrument , för att det internationella valutasystemet skall vara stabilt .
När det gäller argumentet att detta initiativ förstärker osäkerheten är , vad jag förstår , idén med de mycket kortsiktiga kapitaltransaktionerna just att spela på osäkerheten och slå vad om utvecklingen mellan valutor eller mellan olika kortsiktiga ekonomiska tillgångar .
Detta argument förefaller mig därför inte relevant .
Jag skall inte ytterligare gå in på sakfrågan .
Jag tror att alla har sina argument .
Jag vill emellertid fästa er uppmärksamhet på inte bara punkt 9 i resolutionen , utan också punkt 10 .
Vi förväntar oss ett tydligt politiskt ställningstagande med en mycket tydlig tidsfrist , nämligen förberedelserna av höstsammanträdet i Internationella valutafonden , och vi kräver därför , om resolutionen röstas igenom i morgon i kammaren , att kommissionen och rådet kommer till parlamentet och berättar vilka ståndpunkter de tänker försvara vid detta tillfälle .
Fru talman , kära kolleger !
Min grupp gläds verkligen åt att denna debatt äger rum i dag , särskilt som vi inte sparat på ansträngningarna för att tillsammans med kolleger i de olika grupperna uppnå detta .
Vi har naturligtvis inte samma synsätt , och jag tror att vår debatt och de resolutionsförslag vi lagt fram vittnar om det .
Men vi är ändå inte okänsliga för det framsteg som utgörs av kompromissresolutionen , där kommissionen uppmanas att lägga fram en rapport inom sex månader .
Vi tror att Europaparlamentet på detta sätt kan spela sin roll genom att ta initiativet , trots att det är blygsamt , i denna fråga , även om det är självklart - och jag instämmer med föregående talare - att om punkt 9 ifrågasattes , skulle resolutionen naturligtvis förlora hela sitt innehåll .
Vår debatt gäller faktiskt en vital fråga som allt fler medborgare ställer sig på ett berättigat sätt : vilken plats skall vi ge människan och finansvärlden i dagens ekonomi ? 1 800 miljarder dollar , det är värdet av den valuta som varje dag passerar världens växelmarknader , vilket motsvarar mer än en fjärdedel av den årliga världsvolymen av verklig handel med varor och tjänster .
Genom att låta finansen inta en ledande ställning har man ökat kraven på lönsamhet och överallt gjort det svårare att bedriva rörelse .
Det är framtidsperspektivet i det ökande antalet sammanslagningar , förvärv och omstruktureringar av företag , och för de enorma resurserna på finansmarknaderna som bara ökar .
Arbetslösheten och trycket på de anställda i hela världen blir bara värre .
Verklig avsättning och tillväxt förhindras .
Och tillförseln eller det brutala bortdragandet av spekulativt kapital hotar ekonomin i ett stort antal länder , ända till att de faller sönder , såsom i Asien , Ryssland eller Brasilien .
Inför denna nyliberala internationalisering , under finansmarknadernas dominans , ökar kravet , som vår begäran vittnar om , på en annan världsuppfattning där den gemensamma lagen skulle vara skyldighet till solidaritet i en värld där vi blir alltmer beroende av varandra .
Ingen kan bortse från den utmaning för civilisationen som bristen på nära en miljard arbetstillfällen innebär .
Eller behovet av ansträngningar utan motstycke när det gäller utveckling och tillgång till kunskap .
I det hänseendet förtjänar alla idéer att granskas och vi anser att idén om Tobinskatten är en viktig sådan , liksom andra former av tänkbara transaktioner .
Denna skatt kan bidra till att bromsa spekulationen , utan att skada verksamheten i den verkliga ekonomin , och göra det möjligt att lösgöra nya resurser för mänskliga investeringar , i en tid när UNDP uppskattar att det krävs 40 miljarder dollar per år för att utrota fattigdomen , ge alla tillgång till dricksvatten samt tillgodose sanitära behov .
Medan debatten inletts på världsnivå om politikens möjlighet att påverka det ekonomiska området skulle inrättandet av denna skatt kunna bli en av symbolerna för den politiska viljan till att återerövra demokratiska områden som internationella finansaktörer lagt beslag på .
Och jag vill gärna svara kommissionären , som sade att det behövdes ett minimiantal av industriländer för att lyckas med det .
Jag anser att Europeiska unionen består av ett stort antal industriländer och jag tror , liksom Harlem Désir och flera andra talare , att den europeiska union vi utgör kan ta initiativet i det hänseendet .
I vilket fall som helst tror jag att Europaparlamentet skulle berömma sig av att upprepa medborgarnas önskan att kontrollera världen i riktning mot välbefinnande för alla .
Fru talman !
Också jag gläds åt denna debatt som bara dröjt alltför länge .
Vi vet mycket väl att varje generation genom tiderna blint hemfallit åt vad som skulle kunna kallas en dominerande ideologi , dvs. en samling förutfattade meningar som accepteras av den omgivande konformismen , och som ändå till slut visar de kommande generationerna i vilken utsträckning de varit fyllda av dramatiska händelser .
Frihandeln och den permanenta saligförklaringen av internationaliseringen utgör i våra ögon den dominerande ideologin i dag , dvs. det stora misstaget i slutet av vårt århundrade , och är lika farlig som tidigare ideologin med proletariatets diktatur i Kremls korridorer eller , ännu tidigare , den till sanning upphöjda övertygelsen om att jorden är rund .
Vår värld domineras i dag av en enda logik , en enda gud tänkte jag säga , nämligen pengarna i arbete och inte människan i arbete .
Med ett belopp för handel med varor och tjänster som uppgår till 36 000 miljarder francs , dvs. produkten av endast fyra dagars spekulation , har människans producerande verksamhet inte mycket att tacka finansbubblan för .
Den är självförsörjande i ett överbud som överallt fortsätter att förneka människans humanitet , de rikas såväl som de fattigas , även om det är de senare som i slutänden blir uteslutna från de flesta beslutssammanhang , vilka en ytterst liten minoritet lägger beslag på , något som Jean-Pierre Chevènement mycket träffande nyligen kallade " den internationaliserade eliten " .
Det var naturligt att denna elit utesluter all politisk oro från sitt verksamhetsområde och på så sätt kommer undan minsta demokratiska kontroll och i stället helt enkelt lyckas bli både olagliga och oansvariga .
Men folken står emot , vilket deras reaktioner vid det obeskrivliga toppmötet i Seattle vittnar om , där världens ansvariga servilt kom skyndande - med Europeiska kommissionen i täten , tyvärr - och hoppades att deras foglighet vid fötterna av världens härskare Clinton skulle vara tillräcklig för att garantera dem en liten del av kakan .
Utan att räkna med den hälsosamma reaktionen från dem utan rang - individer eller stater - en reaktion som för övrigt var mer organiserad än man sagt , bl.a. i Frankrike tack vare det fantastiska ATTAC-nätet , som kämpar och får allt större genomslagskraft när det gäller att begränsa frihandeln i allmänhet och beskatta internationella finanstransaktioner i synnerhet .
Inrättandet av denna skatt av Tobintyp eller professor Laurés mer realistiska typ , skulle vara politiskt opportun , åtminstone genom sin symboliska betydelse , även om den är låg , eftersom den framför allt skulle betyda att politiken på nytt stabiliseras på ett område som den har uteslutits från , av operatörer vars vinster står i proportion till staternas grad av frånträdande .
Fru talman !
Trots att en del av syftena med Tobinskatten är väl värda att stödjas skulle ett införande av skatten , om detta först i världen och endast sker i Europeiska unionen , innebära en dödsstöt mot den europeiska valutamarknaden .
Om de andra betydande valutahandelsområdena i världen lät bli att införa Tobinskatten , skulle beskattningen i Europa leda till att valutahandeln flyttas över till dessa områden .
Detta har redan klargjorts ett antal gånger under den här debatten .
Det räcker inte med att alla världens industriländer ansluter sig , för då skulle valutahandeln flyttas över till skatteoaser utanför dessa industriländer .
Därför borde ett införande ske globalt .
Det räcker inte med att G7-länderna eller andra industriländer är med .
Att införa skatten både samtidigt och globalt är å ena sidan en så oerhört svår uppgift - och jag personligen tror åtminstone inte att man härvidlag uppnår några resultat - att det vore lika bra att begrava drömmen om införandet av Tobinskatten .
Dessutom , även om man uppnådde enighet om införandet , återstår frågan om uppdelningen av skatteintäkterna .
Centra för valutahandeln i världen kommer knappast att gå med på att skatteintäkterna till exempel via FN används till all världens goda ändamål utan att en betydande andel av skatteintäkterna stannar kvar hos dem .
Vad beträffar möjligheten att genom Tobinskatten förebygga kommande valutakriser måste man lägga märke till att man genom skatten inte avskaffar orsakerna till övervärdering av valutor .
Därför bör man också koncentrera sig på politik - Karas talade också om detta - som leder till att en viss valuta övervärderas i förhållande till sin verkliga potential .
Detta skulle å andra sidan förutsätta en reglering av exporten och importen av kapital , annars skulle det inte vara möjligt att på detta sätt koncentrera sig på politiken .
Trots att Tobinskatten är till synes vettig är den alltså inte problemfri även om man skulle uppnå en överenskommelse om dess genomförande , vilket jag alltså inte tror på .
Man måste komma ihåg att pengar i dag i första hand handlar om information , och att det är kunskapen och det intellektuella kapitalet som i framtiden i allt högre grad kommer att hålla världsekonomin i gång .
Det är därför som de väldiga mängder av kapital som oupphörligen strömmar mellan världens finanscentra inte enbart härrör från spekulativ verksamhet som inte har någonting med den egentliga realekonomin att göra .
Om man med hjälp av sådana arrangemang som Tobinskatt försvårar den här feed back-mekanismens funktion , som alltså ger användarna en möjlighet att välja , kan detta resultera i felaktiga lösningar vars ekonomiska konsekvenser blir så kostsamma att man med hjälp av själva skatten aldrig kan skaffa så mycket .
Därför motsätter sig vår grupp absolut , såsom Karas redan förtjänstfullt konstaterat , att Tobinskatten införs .
Fru talman !
Jag är för beskattning av spekulativa kapitalrörelser över statsgränserna .
Jag tycker att det är alldeles uppenbart att man måste vidta vissa åtgärder .
Under de senaste 30 åren har volymen på valutatransaktionerna blivit 83 gånger större : För det första uppgår alla centralbankers globala reserver knappt till en enda dags valutahandel ; för det andra motsvarar den årliga globala handeln med varor och tjänster bara tre och en halv dagars valutahandel av 350 , dvs .
1 procent av kapitalrörelserna har samband med handel i varor och tjänster och 99 procent är ren spekulation .
De globala valutamarknadernas volym , oförutsägbarhet och irrationella beteende har gjort det svårare och svårare att styra de nationella och regionala ekonomierna .
Datakontrollerade säljprogram som sätts i gång på måfå sätter i gång en lavin som begraver jobb , människoliv och företag över hela världen .
De enda argumenten emot detta är : För det första skulle det försämra valutamarknadens effektivitet - litet besynnerligt med tanke på de profithungriga vansinnigheter vi sett på finansmarknaderna som krossat arbetstillfällen över hela världen : i Östasien , Europa och Latinamerika .
President Chirac har beskrivit de som sysslar med detta som ett aidsvirus i världsekonomin .
Det är nödvändigt att kasta litet grus i maskineriet hos valutaspekulanterna , börsmäklarna och optionshandlarna .
Detta kan naturligtvis inte bara ske i ett land ; det kan inte bara ske inom euroområdet , utan det måste ske på internationell nivå genom globalt samarbete .
Europeiska unionen , Japan och Förenta staterna - euron , yenen och dollarn , skulle kunna utgöra ett sådant block , enligt min mening .
Jag är besviken på EPP-gruppen .
Jag trodde åtminstone att de läste de resolutioner som de röstar om .
Jag är alltså för införandet av en dylik skatt , men det är inte detta omröstningen handlar om i morgon .
Omröstningen i morgon handlar om att vi skall uppmana kommissionen att granska frågan , att undersöka vilka åtgärder och vilka villkor som är nödvändiga i samband med införandet av en dylik skatt .
Jag kan också förstå att kommissionären inte kan stödja en dylik skatt , men jag kan inte förstå varför han inte hade modet att ta tillfället i akt och redovisa sin ståndpunkt genom en granskning av frågan .
Det finns inget som är lika slutet som ett slutet sinne .
Skatten stöds av 47 procent av befolkningen i Förenade kungariket , enligt en nyligen genomförd undersökning av War on Want .
Fransmännen har gett den ett enormt stöd , i synnerhet om den kopplas till ett krav att använda vinsten till att hjälpa utvecklingsländerna med deras ekonomiska skulder och fattigdom .
Parlamentet , rådet eller kommissionen kan inte längre bortse från denna fråga .
Många röster hos folkopinionen kräver nu ett mer genomtänkt svar än : " Det har inte gjorts förut " .
Under det nya millenniet , med nya globala problem som kräver nya globala lösningar , måste de redovisa övertygande skäl till varför det inte går att genomföra nu , i stället för att säga att det inte har gjorts förut .
Fru talman , herr kommissionär , kära kolleger !
En politisk kompromissresolution om nyttan av en skatt på internationella finansiella flöden skulle vara ett första steg mot den nödvändiga trimningen av ett stort antal av våra internationella regler .
Jag har två eller tre punkter jag vill erinra om här .
Ett av huvudkraven från demonstranterna i Seattle var just att inrätta denna typ av skatt , och det är ingen tillfällighet .
Dagens förslag är en stark signal från de rika europeiska länderna som bevisar att de är beredda att avstå från sin egoism , herr kommissionär .
I allas ögon är en sådan solidarisk skatt en rättskaffens åtgärd som inte förhindrar handeln , utan gäller spekulationen och dess snedvridna effekter , kära kolleger till höger .
Detta symboliserar behovet av solidaritet med länderna i söder , särskilt länderna i Afrika , Karibien och Stilla havsområdet som också i stor utsträckning vände sig till oss i Seattle i denna fråga .
För att fullständigt nå sitt mål måste omfördelningen av den valuta som frigörs genom en sådan skatt absolut gå till de fattigaste länderna .
På det viset ger vi ett innehåll dels åt moraliseringen av handelsreglerna dels åt solidariteten med länderna i söder .
Fru talman !
Man kan inte bara ständigt på nytt upprepa antalet , som många av de föregående talarna har gjort , utan man bör också , herr kommissionär , nämna att 80 procent av denna dagliga valutahandel av enorma proportioner inte ligger placerade längre än åtta dagar .
Det kan ju inte fortsätta som i dag att det är mindre lönsamt att investera och skapa arbetstillfällen än att bedriva kortsiktig valuta- och aktiehandel .
Det kan inte fortsätta så att vi förstör de politiska gestaltningsmöjligheter vi faktiskt har .
Det kan inte fortsätta att inkomsterna från icke-ekonomisk verksamhet stiger allt snabbare .
I Tyskland har det , sedan Tobin utvecklade sin idé , visat sig att inkomster från penningtillgångar i dag , utifrån en siffra på 7,6 procent , nästan har fördubblat sin andel av den totala samhälleliga inkomsten .
Det kan ju inte fortsätta så att de fattigaste länderna på jorden är de som utsätts mest för spekulativa påfrestningar till följd av kortsiktiga valutafluktuationer .
Jag tror inte heller att det är ogörligt .
Varför skulle det inte vara möjligt att få till stånd ett avtal mellan G7-staterna , övriga EU-stater , Kina , Singapore och Schweiz angående införande av Tobinskatten ?
Det måste finnas ett allmänt ekonomiskt intresse .
Varför skulle det inte vara görligt att beskatta transaktionerna i valutahandeln med spottar och derivat - alltså de så kallade kassaaffärerna , valutatermin- och optionsaffärerna - särskilt som det är möjligt att utforma ett differentierat system ?
Varför skulle det inte vara görligt att sätta skattesatserna så högt att skatterna inte hotar de på lång sikt ekonomiskt nödvändiga investeringarna och samtidigt slutligen gör de kortfristiga och spekulativa placeringarna oattraktiva ?
Många svåra frågetecken kommer säkert att uppkomma i samband med detta , men det enda riktigt stora problemet hittills som jag kan se är bristen på politisk vilja samt den egoismens princip som visat sig också i dag och består i att skjuta ansvaret ifrån sig på någon annan .
Fru talman !
Vi vill inte ha mer byråkrati , som Karas sade för några minuter sedan .
Vi vill ha lösningar .
Naturligtvis fordrar kapitalmarknaderna tydlighet - det är det som är själva idén .
Tobinskatten kommer att resultera i att det blir öppenhet på ett mycket grumligt område .
" I takt med handelns avreglering , kommer det att krävas fler och fler bestämmelser " , som kommissionär Lamy sade under millennierundan i Seattle .
Han insåg att den inre marknadens och den gemensamma valutans kombinerade effekter , vilka karakteriserar skapandet av Europeiska unionen , är nära förbundna med en enorm mängd nya bestämmelser .
Nu när det är lätt att få tillgång till finansiering över nationsgränserna , är det tydligt att samma förhållningssätt kommer att bli nödvändigt ; i ännu högre grad när vi beaktar att det varje dag omsätts enorma belopp i spekulativt syfte .
Vi världsmedborgare kan inte tillåta den nuvarande spekulationsnivån .
En fortsättning skulle leda till ekonomiskt självmord .
Damer och herrar ledamöter , herr kommissionär !
Man hör ofta att Europa har lyckats uppnå stabilitet i den finansiella sektorn , något som är sant bara om vi begränsar oss till den offentliga sektorn .
Om vi inkluderar även den privata sektorn , kommer vi att märka att vi inte bara har lyckats uppnå denna berömda financial stability , utan att vi också med största sannolikhet sitter på en vulkan som hotar att när som helst få ett utbrott .
Den alltför höga skuldsättningen i den privata sektorn och den motsvarande överdrivna aktieuppgången , de två främsta indikatorerna för stabiliteten på värdepappersmarknaden , har sedan en tid tillbaka kommit in på farligt område , vilket också visas i kommissionens rapport om det ekonomiska läget i Europa , på ett sätt som inte tillåter några tvivel .
Det faktum att allmänheten godtar dessa kurser och inte i panik överger de finansiella marknaderna , kan förklaras med överoptimistiska förväntningar om framtida vinster .
Den spekulativa verksamheten utvecklas bortom all vett och sans och genererar i sin tur vinster , som helt plötsligt kommer att visa sig vara skenbara .
Överoptimismen kommer att ersättas av besvikelse och rädsla , med en börskris , och eventuellt en ekonomisk kris , som följd .
Faran är alltför stor för att vi skall kunna ignorera den .
Vi måste angripa den , hur svårt det än verkar .
Den moderna ekonomiska forskningen har med Tobins och med andras förslag gett oss ett utmärkt instrument , som vi skulle kunna använda oss av , om vi hade den politiska viljan att utarbeta någon slags princip .
Det saknar vi , herr kommissionär .
Den politiska viljan att utforma en princip för att angripa spekulationen .
Den omåttliga dyrkan av eller blinda tron på marknadskrafterna , som liberalerna propagerar för - och jag beklagar att Gasòliba i Böhm har gått - , kan inte fortsätta att i all evighet styra demokratin , för den styr den rakt mot katastrofen !
Fru talman , herr Bolkestein !
Det är faktiskt rent utsagt otroligt vilken okunnighet man diskuterar med här .
Vi behöver en grekisk kollega för att någon äntligen skall säga vad den här Tobinskatten egentligen handlar om .
Ni avslår den utan vidare eftersom ni inte förstår någonting av det .
Att högern är emot skatter är självklart , men de skulle aldrig ha fått överföra dessa miljon- och miljardbelopp till Schweiz .
Det är självklart !
Nu uppmanar jag er , helt medvetet , att lämna ett bidrag för att stoppa det spekulativa finanskapitalet och äntligen motarbeta long term projects med hjälp av long term capital .
Det har aldrig gjorts i Sydostasien och det har aldrig gjorts i Europa , och att kollegan Karas från Österrike inte längre är här förstår jag också med tanke på deras finansiella agerande .
Det är samma gamla skit !
Vi behöver en Tobinskatt , så att vi kan ingripa med skatteinstrumentet !
Fru talman , jag är oerhört sur över kommissionens politiska okunnighet , dvs .
Bolkesteins politiska okunnighet !
Med den inställning han har till Tobinskatten borde han fundera på varför han överhuvudtaget är här !
Fru talman !
Jag har också delvis upplevt debatten som riktigt skrämmande .
Det kanske inte är en slump att det inte finns någon kvar av de konservativa , för det man företrätt under beteckningen marknadsfrihet har inte längre någonting att göra med de respektingivande principerna för den sociala marknadsekonomin , som skänkt oss ett sådant välstånd under gångna årtionden .
Fortsätter vi med att på det här sättet förklara finansmarknaderna för heliga , vilket ideologin säger , ja om vi till och med påstår att varje ingrepp i dessa marknaders funktion är emot framsteg och tillväxt i ekonomin så har vi helt visst slagit in på fel väg , och det kan bli riktigt farligt med tiden .
De som sitter på penningtillgångar samlar för närvarande på sig allt större förmögenheter , vilka i sin tur kräver att bli placerade .
Vi har att göra med en asset inflation av global omfattning .
På så sätt uppstår det ständigt spekulationsblåsor på finansmarknaderna , vilka medför ökad ekonomisk oro som i sin tur utgör en fara för ekonomin i stort .
De som blir lidande av detta är de medelstora företagen och många arbetstagare .
Men det finns botemedel mot detta , det är möjligt att göra något .
Ett minimum för att det skall gå är dock att det görs seriösa studier , inte från kommissionens sida utan också av verkligt ekonomiskt renommerade inrättningar över hela Europa .
Också det är något genomförbart .
Och då skall man inte hela tiden välja fel personer för sina argument .
Att Tobinskatten inte skulle vara tekniskt genomförbar stämmer inte - i datorernas tidsålder går det .
Att skatteoaserna mycket ofta inte är något annat än minnen i maskinvaruform för stora europeiska banker bör man inte heller bortse ifrån .
Sammanfattningsvis : Vi får inte tillåta att realkapital och finanskapital fjärmar sig alltför långt från varandra , annars lär vi på sikt närma oss förhållanden som vi redan upplevt flera gånger på den här kontinenten och som lett till fruktansvärda katastrofer .
( Applåder ) Fru talman , bästa kolleger !
Låt oss beskatta valutaspekulationen , den producerar inte någonting nytt .
Skatten skulle rikta sig mot helt rätt objekt : spekulanterna .
Vem är det som försvarar dessa spekulanter samtidigt som sjuksköterskor och lärare betalar höga skatter ?
Artikel 73 c i Fördraget om Europeiska unionen gör det möjligt att beskatta transaktioner .
Kapitalskattens motståndare stödjer dessa skatteflyktscentraler , skatteparadis , vars antal sammanlagt uppgår till 62 .
Unionen borde skapa ett skatteavtal som vilka länder som helst skulle kunna ansluta sig till i början .
En låg Tobinskatt skulle inte förorsaka några större problem med skatteflykt .
Det är ett märkligt påstående att man inte kan skapa en skatt om inte alla ansluter sig .
Det var också bara några få stater som grundade Europeiska unionen , och ni ser hur det ser ut i dag .
Faktum är att det största problemet är politiskt - man vill inte beskatta kapitalet utan skärpa beskattningen av människorna .
Skatten skulle slutgiltigt politisera det globala , odemokratiska finansmaktssystemet .
Vi måste , bästa kolleger , utmana världens spekulationselit , som med ensamrätt vill leda världens ekonomiska planering genom att hålla sig utanför skattesystemen . .
( NL ) Fru talman !
Får jag till att börja med tacka alla talare och allra först naturligtvis Désir så innerligt för att den här debatten äger rum i kväll .
Vad man än må tänka om samtalsämnet så är det tydligt att det är ett viktigt ämne .
Det är också därför som det varit på tapeten i flera år nu och det är tillfredsställande att kommissionen i kväll kan ge ett svar på det här .
Jag skulle vilja börja med att ta upp två anmärkningar från parlamentsledamoten Gasòliba .
Han har sagt att globalisering är ett positivt fenomen och det håller jag med honom om .
Jag tror att globaliseringen bidragit till att många länder som hittills stod vid sidan av strömmarna i världshandeln nu deltar i den , nu har blivit en del av världshandelssystemet och så vitt jag vet har inget land någonsin fått det sämre på grund av internationell handel .
Jag ser alltså globaliseringen som något positivt , vilket Gasòliba också sade , och jag anser att den har bidragit till den nya internationella arbetsfördelning som många strävat efter i flera år .
En andra anmärkning från Gasòliba var att det för ögonblicket inte finns några bevis för att Tobinskatten skulle stabilisera valutakurserna .
Det tror jag att han har rätt i .
Jag känner heller inte till något skäl till varför en beskattning av valutakurstransaktioner skulle leda till att de stabiliserades .
Jag tycker att det är två viktiga anmärkningar , det är därför som jag upprepar dem nu .
Vidare skulle jag , fru talman , vilja påpeka att ingen av talarna i kväll har fört fram något samband mellan Tobinskatten å ena sidan och Europeiska unionens funktion å den andra .
Vi känner ju alla till Romfördraget .
Vi vet ju att en av friheterna är fri rörlighet för kapital .
Fru talman !
Jag kan tala om för parlamentet att mitt dagliga arbete bland annat består i att jag tillsammans med mina avdelningar och mina kolleger försöker integrera de finansiella marknaderna i Europa helt och hållet så att den finansiella rörligheten blir så lätt och smidig som möjligt .
I min funktion är jag alltså en motståndare till alla åtgärder som skulle kunna försvåra den finansiella rörligheten .
Då kan ni väl ändå inte förvänta er av den här kommissionären att han skulle instämma med en skatt som skulle innebära just ett hinder för den internationella ekonomiska rörligheten .
Enligt min åsikt strider alltså Tobinskatten mot Romfördraget och det är en viktig teoretisk invändning som ingen av talarna tagit upp i kväll .
Fru talman !
Efter dessa , tycker jag , ganska grundläggande anmärkningar finns det också praktiska invändningar mot Tobinskatten och dessa har bland andra Karas tagit upp .
Man har , tyvärr tycker jag , anmärkt att Europeiska unionen internt inte lyckats komma överens om vissa skatteåtgärder .
Det visar hur besvärliga dessa ärenden är .
Om vi inte ens internt har kunnat komma överens hur skall vi då kunna övertyga andra handelspartner ?
Det kommer att bli svårt , tror jag .
Fru talman !
Jonckheer sade att det här skulle kunna vara en åtgärd för stabilisering av de finansiella marknaderna .
Jag tror dock att vi här har att göra med ett symptom och att vi måste undersöka orsakerna , att det är bättre att försöka åtgärda orsakerna än att försöka göra något åt symptomen när det troligen inte heller är möjligt och , som sagt , när det helt säkert strider mot Romfördraget .
För att få bort de här orsakerna måste man se efter vad som händer i de berörda länderna .
Är det så att de länderna kan prunka med vad man på engelska kallar för good governance ?
Är det så att räntan är låg och inflationen är låg ?
Att marknaderna för produktionsfaktorer , bland annat arbetsmarknaden , fungerar smidigt ?
Det är inte alltid fallet .
Vill vi alltså undersöka orsakerna till de instabila valutakurserna så måste vi kunna se beståndsdelarna i en good governance och rikta vår första uppmärksamhet mot dessa .
Dessutom , och det har också redan tagits upp av till exempel Gasòliba I Böhm , men också av andra , behövs det mer kontroll .
Mer nationell kontroll , nationella regeringars kontroll av nationalbanker och även internationellt , till exempel genom Internationella valutafonden ( IMF ) .
Jag tror alltså att vi bäst tar oss an orsakerna genom att å ena sidan se till att det i de berörda länderna förs en good governance och å andra sidan att det kommer mer nationell och internationell kontroll för att undvika sådana urspårningar .
Olika parlamentsledamöter har sagt att det ändå måste anslås mer pengar för stora projekt .
Kreissl-Dörfler talade till exempel på engelska om long term financing for long term projects - det är en självklar fråga .
Mitt svar är att länderna i första hand borde göra vad de lovat att göra , nämligen anslå 0,7 procent av sin bruttonationalprodukt till bistånd och utvecklingssamarbete , så att mycket mer pengar än nu kan användas för sådana long term-projekt via den väg som är bestämd för det ändamålet , nämligen bidrag till utvecklingssamarbete och inte via en konstgjord och troligen skadlig väg , nämligen Tobinskatten .
Fru talman !
Jag skulle gärna vilja sluta där .
När det gäller den resolution som jag sett ett utkast till så avvaktar kommissionen omröstningen och skall på grundval av den bestämma sin ståndpunkt och jag tackar er för tillfället att delta i den här debatten .
Jag har mottagit fyra resolutionsförslag , som inlämnats på grundval av artikel 40.5 i arbetsordningen .
Fru talman , dessvärre är jag inte lika bra som ni på franska .
Det skulle dock glädja mig om Bolkestein kunde lyssna helt kort , vilket inte verkar vara möjligt eftersom han just nu talar med Randzio-Plath .
Kan ni göra honom uppmärksam på att jag vill säga en sak till honom ?
Monsieur Bolkestein , je veux vous dire quelque chose !
Dessvärre är jag inte lika bra på nederländska som ni .
Men jag skulle ändå vilja säga er något .
Det är faktiskt inte fråga om ett initiativ bara för att irritera kommissionen , detta att vi är för en Tobinskatt .
Vi vill undersöka möjligheterna att införa en Tobinskatt .
Det skulle bara vara ett bland många andra instrument .
Förhoppningsvis finner vi också er på vår sida när det gäller detta .
Politiskt sett har jag alltid svårt för när folk säger att det behöver vi inte , det vill vi inte och det kan vi inte .
Det är inte er uppgift att bestämma det , utan vår .
Vilket också hänger samman med den nyväckta självkänslan hos parlamentet .
Om det skulle jag gärna diskutera med er , varken mer eller mindre .
Vi kan strunta i alla andra utsvävningar , men jag respekterar er som seriöst sinnad kommissionär som vill ta sitt arbete på allvar .
Men respektera då också oss som ledamöter som vill ta vårt arbete på allvar , och till detta hör Tobinskatten !
Fru talman !
Det verkar föreligga ett förbiseende och i förteckningen över inlämnade resolutionsförslag som ni just nämnt ingick inte det gemensamma förslaget till kompromissresolution från PSE-gruppen , den liberala gruppen , GUE-gruppen , Gruppen De gröna samt Kuntz och Coûteux .
Kära kollega !
Jag noterar ert uttalande och förekomsten av denna gemensamma resolution .
Om ordförandeskapets enheter bekräftar att den lämnats in , skall den självfallet beaktas .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum på torsdag kl .
12.00 ( Sammanträdet avslutades kl .
20.14 )
