 
Återupptagande av sessionen Jag förklarar Europaparlamentets session återupptagen efter avbrottet den 21 januari 2000 .
Fru talman !
Tillåt mig påminna om att i morgon är det två år sedan katastrofen i Cermis .
För två år sedan kapade ett amerikanskt flygplan från Natobasen i Aviano under en övningsflygning på låg höjd - under den tillåtna säkerhetsgränsen - linorna till en linbana i Cavalese i Italien och orsakade över 20 europeiska medborgares död .
Alltsedan dess väntar offrens familjer , som inte har kunnat söka tröst i någon rättvisa eftersom den ansvarige piloten inte har fått något straff , på att få åtminstone ekonomisk ersättning från USA .
Jag vill därför uppmana parlamentets talman och rådets ordförande att hos de amerikanska myndigheterna utverka en omedelbar ersättning i enlighet med de rättigheter som offrens familjer har .
Tack , fru Angelilli !
Jag noterar ert inlägg .
 
Föredragningslista Nästa punkt på föredragningslistan är fastställande av arbetsplanen .
Efter den begäran jag erhållit från flera politiska grupper och efter den talmanskonferens vi just haft , föreslår jag en debatt på en och en halv timme om en aktuell och brådskande fråga av större vikt , i enlighet med artikel 50 i arbetsordningen , om unionens reaktion på regeringsförhandlingarna i Österrike .
Om ni beslutar att föra upp denna debatt på föredragningslistan kommer den att inledas av rådets ordförande Seixas da Costa och kommissionens ordförande Romano Prodi .
Vill någon uttala sig för detta förslag ?
Fru talman !
Jag vill göra ett inlägg för att uttala vårt stöd för talmanskonferensens beslut , och med tanke på att jag kritiserade ordförandeskapet offentligt i januari , ta tillfället i akt för att tala om att jag i dag , personligen och som företrädare för Europeiska socialdemokratiska partiets grupp , anser att ordförandeskapet har gjort högst adekvata uttalanden i denna fråga , och att vi i alla avseenden är eniga i dessa .
( Applåder ) Mot bakgrund av detta , fru talman , är det svårt att tänka sig en debatt som bättre överensstämmer med det som står i artikel 50 i parlamentets arbetsordning .
Detta är en aktuell debatt , som är oerhört viktig och brådskande .
Vi anser därför att den bör tas med på föredragningslistan .
( Applåder ) Finns det någon kollega som vill uttala sig emot detta förslag ?
Fru talman !
Jag vill uttala mig emot av principskäl som förefaller mig fullständigt grundläggande , eftersom det handlar om att respektera fördragen , bl.a. artikel 7 i Amsterdamfördraget .
Fru talman , kära kolleger !
Vi har hittills trott att Europeiska unionen , enligt bestämmelserna i Rom- och Parisfördragen genom vilka gemenskaperna grundades , och som sedan blev unionen , var en sammanslutning av fria , oberoende och suveräna stater .
Även om ett stort antal förändringar gjorde att vi betvivlade detta , har vi ändå ansett att detta var fallet och nyligen hänvisade man återigen till subsidiaritetsprincipen , även om det var halvhjärtat .
Fru talman !
Det förefaller emellertid i dag uppenbart att om man inleder den debatt som ni och talmanskonferensen ber oss att inleda , på grundval av artikel 50 , skjuter man en fruktansvärd bräsch i principen om frihet , staternas suveränitet och regeringarnas fria sammansättning , som är resultatet av demokratiska val , och då kan i morgon en annan majoritet i parlamentet lägga sig i bildandet av en regering som ändå är resultatet av fria , regelrätta , fredliga och demokratiska val inom en medlemsstat .
Om ni ratificerar ...
Herr Gollnisch !
Ursäkta mig , men ni har bara en minut .
Jag vet att ni alltid är noga med att arbetsordningen skall respekteras .
Fru talman !
Jag trodde att jag hade tre minuter .
Jag ber om ursäkt .
Om ni ratificerar denna utveckling ratificerar ni utvecklingen av en union i riktning mot en organisation som kommer att bryta mot suveräniteten och friheten för medlemsstaternas nationer , och vi har då inget annat val än att utträda ur en sådan union .
Vi har lyssnat till en talare för och en talare emot .
Jag kommer nu att låta förslaget till ändring av föredragningslistan gå till omröstning .
( Parlamentet biföll begäran . )
( Applåder ) Debatten har placerats i början av föredragningslistan .
 
DEBATT OM AKTUELLA OCH BRÅDSKANDE FRÅGOR Nästa punkt på föredragningslistan är den aktuella och brådskande debatten om frågor av större vikt .
 
Regeringsförhandlingar i Österrike Nästa punkt på föredragningslistan är debatten om regeringsförhandlingarna i Österrike .
Jag ger genast ordet till rådets ordförande .
Fru talman , ärade kollegor !
Av Europeiska unionens portugisiska ordförandeskap har jag blivit ombedd att tillsammans med parlamentet uttala vår mening rörande det politiska läget i Österrike och vilka konsekvenser detta har för förbindelserna med de övriga unionsländerna .
Först och främst vill jag klargöra att när det gäller den portugisiska premiärministerns uttalande den 31 januari , som företrädare för tre andra länder som också är unionsmedlemmar , så är det fråga om en gemensam politisk ståndpunkt antagen av fjorton stats- och regeringschefer företrädda av Portugal .
Texten i den gemensamma ståndpunkten är väl avgränsad med ett klart och tydligt syfte : den bilaterala förbindelserna mellan de fjorton länderna och en österrikisk regering som delvis kommer att bestå av landets liberala parti .
Jag vill påminna om vad som då sades .
1 - De fjorton medlemsstaternas regeringar kommer varken att främja eller acceptera officiella bilaterala förbindelser på politisk nivå med en österrikisk regering där Österrikiska liberala partiet ( FPÖ ) ingår .
2 - De österrikare som sitter på poster i internationella organisationer kan inte räkna med något stöd från de fjorton länderna .
3 - De österrikiska ambassadörerna i unionens huvudstäder kommer enbart att tas emot å yrkets vägnar .
Jag tror att man under de senaste dagarna mer än väl har klargjort skälen till de fjorton ländernas gemensamma ståndpunkt .
Först och främst ländernas gemensamma tolkning av den interna politiska situationen i Österrike , där man drog slutsatsen att ett inkluderande av ett parti som FPÖ skulle kunna förändra respekten för de gemensamma värden som unionens medlemsländer har lovat att värna .
Ingen känner till Jörg Haiders officiella ståndpunkt och de mera konkreta politiska idéer som respektive parti försvarar .
Jag tycker det är onödigt att påminna om deras ursäktande inställning till den nazistiska regimen , deras attityd gentemot utlänningar och invandrare och deras framhållande av en populistisk nationalism som påminner om forna dagar .
Vår tolkning är att ett sådant parti har en helt annan ståndpunkt än den som vi förespråkar i Europa och som för övrigt är den som unionen valt att föra fram i sina externa förbindelser , såväl inför den kommande utvidgningen som när det gäller den gemensamma utrikes- och säkerhetspolitiken .
Man kommer att säga att den nuvarande situationen har uppstått på grund av det österrikiska folkets fria val , vilket måste respekteras för att undvika en inblandning i landets interna angelägenheter .
För det första , herr talman , ärade kollegor , ingen ifrågasätter en demokratiskt vald regim i Österrike eller det senaste valresultat .
Valresultatet visar , och det är bra att det kommer fram , att en stor majoritet av österrikarna fortfarande är emot Jörg Haiders parti .
Vad vi menar och beklagar är att man i en sådan situation valt en regeringslösning som sätter delar av landets politiska makt i händerna på ett parti vars ledare inte på något vis värnar om de grundläggande principer Österrike lovat att respektera , värna och främja .
( Applåder ) Österrike har all rätt att välja sin egen regering , men vi har samma rätt , och skyldighet , att säga vår mening om de politiska alternativ som vi menar avviker från de löften Österrike på ett internationellt plan har avlagt .
Detta gäller i dag för Österrike liksom i morgon för vilket annat land som helst inom Europeiska unionen .
( Applåder ) Jag upprepar : Detta gäller i dag för Österrike och i morgon för vilket annat EU-land som helst .
Å andra sidan vet vi alla i dag att frågor om mänskliga rättigheter , de grundläggande rättigheterna , de stora demokratiska principerna samt rättsstaten , minoritetsskyddet och kampen mot rasism , främlingsfientlighet och intolerans inte bara är frågor för de inhemska domstolarna .
I synnerhet när landet i fråga är en del av en statsgemenskap som grundar sig på detta i sitt civiliseringsprojekt .
Det Europa som vi vill bygga och befästa är inte längre bara ett ekonomiskt projekt , utan en gemenskap med värden och principer baserad på en politisk union och ett inrättande av ett stort område för frihet , säkerhet och rättvisa där solidariteten sätts i förgrunden .
( Applåder ) Fru talman , ärade kollegor , därför menar vi att det är såväl vår rättighet som skyldighet att berätta för våra österrikiska vänner , som för övrigt länderna utanför Europeiska unionen har gjort , att deras regeringsval måste få vissa påföljder för våra framtida relationer eftersom Haiders parti fick ingå i deras regering .
Beträffande de konkreta påföljderna , där kommissionens uttalande från i går gav vissa ledtrådar , kommer Europeiska unionen att försöka fortsätta att arbeta och bevara den sanna respekten för fördragen samtidigt som den österrikiska regeringens agerande noggrant kommer att granskas .
Gemenskapen är ett mycket speciellt område , reglerad av synnerligen konkreta rättspolitiska lagar , och måste därför bemötas på ett särskilt sätt .
( Ihållande applåder ) Fru talman , mina damer och herrar !
Kommissionen sammanträdde i går morse och fattade , självständigt och med stöd från samtliga medlemmar i kollegiet , politiska beslut av grundläggande betydelse .
Redan i går förklarade sig kommissionen dela den oro som unionens 14 medlemsstater gav uttryck för och som upprepats här av företrädarna för ordförandeskapet .
I dag , inför er alla , och som företrädare för hela kommissionskollegiet , kan jag upprepa detta .
Låt mig i första hand med kraft rikta er uppmärksamhet på det som i ett ögonblick som detta är kommissionens politiska roll .
På samma sätt som parlamentet , är kommissionen en av unionens övernationella institutioner och kan just därför inte ha några bilaterala diplomatiska förbindelser med medlemsstaterna .
Det är just när kontinuiteten , sammanhållningen och försvaret av unionens gemensamma värderingar verkar hotade , som kommissionens politiska roll upplevs som starkast och tydligast .
Låt oss inte glömma , mina damer och herrar , att Romfördraget inte innehåller någon artikel om utträde , vare sig frivilligt eller påtvingat , för en medlemsstat .
Och skälet till detta är att själva grundtanken med den fantastiska konstruktion som kallas Europeiska unionen är just att varje enskild stat , i det ögonblick som man blir medlem i unionen , fullständigt och för alltid skall acceptera unionens grundläggande principer .
Dessutom beskriver fördragen i detalj vilka åtgärder som skall vidtas för att de principerna verkligen skall respekteras .
Mot den bakgrunden skulle kommissionen frånsäga sig sitt ansvar om den skulle försöka bibehålla arbetsrelationer med Österrike , på samma sätt som med alla de övriga medlemsstaterna .
Mina damer och herrar !
När någon av unionens medlemsstater befinner sig i svårigheter , är det hela unionen som befinner sig i svårigheter .
( Applåder ) Den skyldighet som en stark övernationell institution har är inte att isolera enskilda medlemsstater , utan att oupplösligt binda dem vid unionens grundläggande värderingar .
Den skyldigheten kommer kommissionen att hävda med den yttersta kraft .
Å andra sidan finns det ingen anledning att uppmana kommissionen att fortsätta följa utvecklingen i Österrike , steg för steg .
Europeiska unionen kan inte överleva utan principerna frihet , demokrati och respekt för mänskliga rättigheter .
Det är unionens grundvärderingar .
De är själva unionens existensberättigande , de är frukten och resultatet av de högtidliga löften som medlemsstaterna har avgivit när det gäller att respektera människor och folk , oavsett tro , ursprung eller samhällsställning .
Dessa principer överensstämmer helt med respekten för rättsstatens principer och kommissionen , som är garanten för rättsstaten , kommer inte att vika en tum när det gäller dess försvar .
Även det mest obetydliga intrång när det gäller människors eller någon minoritets rättigheter kommer vi att reagera på med kraft .
Som en ledamot i ett av kandidatländernas parlament sade till mig , så är Europa en union av minoriteter och känner därför en djup respekt för alla enskilda individers rättigheter .
Fru talman , mina damer och herrar !
Tillåt mig ännu en mycket kort reflexion .
Med sina över 900 år är universitetet i Bologna , mitt alma mater , och det äldsta universitetet i världen .
På väggarna i en av de vackraste salarna kan man fortfarande se vapensköldarna från de studenter och lärare som valde det universitetet , för hundratals år sedan , som sitt lärosäte .
Där finns fortfarande över 7000 vapensköldar från hela Europa , från Transsylvanien till England .
Detta var redan då Europa : en plats där idealen inte kände av några av den tidens geografiska och politiska gränser , en gemenskap med gemensamma värderingar , ideal och kunskaper .
Men Europas historia har inte vävts samman enbart av kulturellt utbyte , kunskapens utvidgning och en robust , gemensam värdegrund .
Bredvid vapensköldarna från de olika universitetssamfunden , i varje liten by i Europa , bär monumenten över dem som fallit i kriget vittne om de tragedier som drabbat vår kontinent .
Europas historia har under sekler utmärkts av en obruten följd av krig och konflikter .
Europa , civilisationens vagga , har gjort sig skyldigt till de mest avskyvärda missdåd som förekommit i mänsklighetens historia .
Därför valde jag att som första handling under mitt ordförandeskap göra en pilgrimsfärd till Auschwitz , för att klart och tydligt , men ändå med den stillhet som platsen kräver , påminna om att detta är minnesplatsen framför alla andra , att Europa inte får glömma , och för att upprepa att dagens och morgondagens Europa är , och inte någonsin kommer att kunna vara annat än , en union av frihet , rättvisa , säkerhet och fred .
Frihet , rättvisa , säkerhet och fred .
Detta är vad Europeiska unionen har varit och det som Europeiska unionen förblir .
Den mest enastående , modiga och framgångsrika politiska konstruktionen under det sekel som just har avslutats har kunnat garantera sina medborgare frihet , rättvisa , säkerhet och fred .
Och det är detta som ett enat Europa vill erbjuda under det sekel som just har inletts , till dem som förbereder sig för att vara en del av det .
I dag på eftermiddagen , just i detta ögonblick , borde jag egentligen ha befunnit mig i universitetet i Lovanio för att tillsammans med den franske premiärministern och generaldirektören för Världshälsoorganisationen , fru Brundtland , promoveras till hedersdoktor .
Jag kommer att komma litet för sent till den ceremonin , men jag tror att det inte finns ett bättre sätt att hedra ett universitet , som är en av den europeiska kunskapens mest betydelsefulla symboler , än att komma hit , till detta parlament , det högsta uttrycket för folkligt självbestämmande , och vittna om detta passionerade engagemang , mitt personliga och Europeiska kommissionens , när det gäller försvaret av de principer som utgör själva grunden för ett enat Europa .
( Applåder ) Fru talman , herr kommissionsordförande , herr rådsordförande , kolleger !
Europeiska folkpartiets grupp ( kristdemokraterna ) och Europademokraterna följer händelserna och diskussionen om utvecklingen i Österrike med oro och spänning .
Vi har i vår grupp - det erkänner jag gärna och jag anser att det är ett tecken på styrkan i vår grupp - fört en lidelsefull debatt , och aldrig har det i samband med ett problem eller ett ärende begärts ordet så många gånger som i dag i vår grupp , och jag tackar alla kolleger som har yttrat sig så seriöst .
En sak bör stå klart : Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater är ense i sin kritik av flera uttalanden från FPÖ : s ordförande i Österrike .
Vi fördömer hans taktlöshet de senaste dagarna , i synnerhet gentemot den franske presidenten Jacques Chirac och den belgiska regeringen .
Vi tillbakavisar detta med all bestämdhet !
( Applåder ) Vi , PPE-DE-gruppen , försvarar människornas värdighet , rättsstaten , demokratin och friheten , och dessa principer och värderingar försvarar vi mot ytterligheter både åt höger och vänster .
( Applåder ) Kristdemokraterna , som är en viktig kärna i vår grupp - och detta är det kanske inte många som känner till - uppstod ur motståndet mot nationalsocialismens totalitära system , som också var människoföraktande , men även mot det totalitära systemet hos den människoföraktande kommunismen .
( Applåder ) Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater företräder också i dag de värderingar som hystes av dem som lade grunden till Europas enande - Robert Schuman , Alcide de Gasperi , Konrad Adenauer och Winston Churchill , och det fanns många flera - och dessa värderingar , som fanns bland dem som grundlade Europa , är våra värderingar även år 2000 .
Dessa principer utgör också måttstocken för de bedömningar som vi gör i fråga om aktiviteterna och agerandet och orden i medlemsstaterna och även hos våra regeringar .
Här vill jag säga : Vi har förtroende för våra österrikiska vänner i det österrikiska europeiska folkpartiet .
( Applåder ) Man måste påminna om att det österrikiska folkpartiet mer än något annat parti under Alois Mock och Wolfgang Schüssel - den ene var ekonomiminister och den andra utrikesminister - har berett väg för Österrike in i Europeiska unionen .
Vi minns att år 1998 , och det är ju inte länge sedan , yttrade sig alla här i parlamentet positivt om Österrikes ordförandeskap , och Wolfgang Schüssel , ordföranden i ÖVP ( Österrikiska folkpartiet ) agerade här särskilt lidelsefullt och engagerat .
Nu har Österrike haft val , och jag anser att det inte är någon mening med att skälla på väljarna .
Man måste också erinra om att det ju förts förhandlingar med SPÖ ( Österrikiska socialdemokratiska partiet ) .
Jag beklagar att dessa inte var framgångsrika , men varför var de inte det ?
Eftersom den del av SPÖ som var fackföreningsorienterad inte var beredd att stödja det som förbundskansler Klima hade garanterat ...
( Applåder från höger , högljudda tillrop från vänster ) ... , nämligen ett saneringsprogram för ekonomi och finanser .
Detta är sanningen , och hur högljutt ni än ropar , så kan ni inte sopa detta under mattan med hjälp av missnöjesyttringar !
Vi förväntar oss att en regering under ÖVP : s ledning , om det blir så , företräder och genomför de värderingar och principer som Europeiska folkpartiet har , och dessa principer är ett otvetydigt erkännande av alla människors värdighet och en uppmaning till tolerans gentemot alla människor , och i synnerhet också en konsekvent fortsättning på politiken att ena Europa , vilket Republiken Österrike på ett föredömligt sätt har gjort i flera årtionden .
Vi kommer att mäta den österrikiska regeringens handlande , om den kommer att ledas av ÖVP , på hur man garanterar rättsstaten , demokratin och friheten , och vi vill uttryckligen tacka er , herr kommissionsordförande och hela kommissionen för att ni inte först i dag avgav ett klokt och balanserat yttrande som motsvarar Europeiska unionens fördrag , utan att ni gjorde det redan i går .
Vi står vid er sida när ni uppfattar er som en väktare av fördragen , och låt oss därför gå denna väg gemensamt !
Det förväntar vi oss och säger som Europeiska folkpartiet grupp ( kristdemokrater ) och Europademokrater : Vi vill ha ett rättens Europa , vi vill ha ett fredens Europa , vi vill ha ett toleransens Europa !
Vi vill inte ha något isolerat Europa , utan vi vill föra samman Europas folk , så att vår kontinent på 2000-talet får en framtid i frihet , demokrati och fred !
( Livliga applåder från PPE-DE-gruppen ) Fru talman , herr kommissionsordförande , herr tjänstgörande rådsordförande !
Europeiska socialdemokratiska partiets grupp vill härmed förmedla tre budskap till den europeiska allmänheten .
Det bör påpekas att vi är helt överens i samtliga tre fall .
För det första vill vi uttala vårt fulla stöd och vår uppbackning av det uttalande som har gjorts av rådets tjänstgörande ordförandeskap och 14 medlemsstater , för vi anser att detta är i linje med den värdegemenskap som vi alla , inte bara en politisk maktfaktor , har skapat .
Hur som helst är det en värdegemenskap som utgör en antites till den som försvaras av det parti som ironiskt nog kallas Österrikiska liberala partiet .
Det Europa som vi är på väg att bygga upp grundar sig på de bittra erfarenheter som vi alla har gjort , och Europeiska socialistiska partiets grupp fördömer de förolämpningar som har lanserats mot den franska republikens president och mot den belgiska regeringen , men även mot socialisterna , för även vi är europeiska medborgare , och i dag , mina damer och herrar , talar man om de österrikiska socialisterna som landsförrädare .
Och en sak vill jag påpeka för er : jag var själv under många år en landsförrädare , åtminstone enligt general Franco .
( Applåder ) Även president Guterres förrådde Salazar , och det tror jag även Europeiska folkpartiets grupp måste medge och hävda .
Dessutom , anser jag att kommissionen , ordförande Prodi , har varit fördragens väktare .
Men jag vill påminna ordförande Prodi om att han i utnämningsdebatten talade om kommissionen som en europeisk regering .
En regering måste vissa större beslutsamhet och större mod .
Det uppmanar jag i dag ordförande Prodi att göra .
( Applåder ) Med all respekt för en sådan kompetent kommissionär som Fischler , skulle jag med tanke på de , språkligt motiverade motsägelsefulla uttalandena angående ordförande Prodis eventuella begäran om Fischlers avgång , uppskatta ett klargörande inför parlamentet i den frågan .
För det andra , fru talman , vill vi framföra ett mycket tydligt budskap till det österrikiska folket .
En uppmaning till den majoritet av den österrikiska befolkningen som inte har röstat för Haider , som har röstat för demokratiska alternativ som innebär att man tar ställning för Europa - och jag måste påpeka att även om Schüssel var finansminister , så bidrog även förbundskansler Vranitzky till Österrikes integrationsprocess .
Man får inte vara så sekteristisk på det politiska området .
Österrikes inträde i gemenskapen är något vi har åstadkommit tillsammans .
Det var allas , inte bara en enskild grupps verk .
Därför , fru talman , anser jag att vi har både en rättighet och en skyldighet att kräva att österrikarna noga överväger och ifrågasätter detta , för en farsot av det slag som vi redan har drabbats av i Europa är inte bara skadlig för Österrike , utan kan även sprida sig och då syftar jag på historien .
Därför skulle jag vilja veta om PPE , förutom sitt försvarstal för Schüssel , som skall ge oss alla garantier , precis som Chamberlain och Daladier i München år 1938 , har tänkt vidta några åtgärder gentemot det österrikiska konservativa partiet om det fortsätter med detta vansinniga projekt .
För det tredje , om vi inte protesterar mot denna förnuftsvidriga allians , kan jag lova , mina damer och herrar , att vi lika gärna kan ge upp Europeiska unionens främsta målsättning , utvidgningen , för vad skulle ni tycka , om ni vore tjecker eller slovener eller ungrare och hade en granne som bemötte er med en rasistisk attityd och inte ville att ni blev medlemmar ?
Därför tror jag , mina damer och herrar , att det här är en viktig dag för det politiska Europas begynnelse .
Vi stöder rådet och anser att det är vår rättighet och skyldighet att vända oss till det österrikiska folket , för att de allvarligt skall överväga detta vansinniga alternativ .
( Applåder från PSE ) Fru talman !
Min grupp välkomnar denna debatt för den är betydelsefull .
Detta är första gången i det moderna europeiska projektets historia som vi börjar se ett parti från extremhögern integreras i politiken .
Det är djupt oroande .
FPÖ hävdar att om man läser deras litteratur och deras programförklaring finns där mycket som man skulle kunna känna sig delaktig i .
Så är det kanske men låt mig i dag föra till protokollet den långa och svåra upplevelse som vi liberaldemokrater genomgick med österrikiska FPÖ inom vår familj Liberal International .
Så tidigt som 1986 hade vi anledning tro att Jörg Haider inte var en man vars principer eller inställning överensstämde med anständighet och modern liberalism .
I november 1991 efter en lång intern debatt inom Liberal International och många besök i Wien för att diskutera frågor avstängde vi temporärt FPÖ som medlem och i juli 1993 uteslöt vi dem .
( Applåder ) Vi uteslöt dem då och vi fortsätter att förkasta det som Haider står för nu .
Låt mig berätta för er vad vi lärde oss under denna långa erfarenhet .
Det fanns många bland oss som sade " läs texten " .
Det fanns många fler bland oss som sade " läs undermeningen " , " se på kontexten " .
Ord som används i politiska sammanhang kan vara uppviglande , kan vara upphetsande eller försonande .
Vi ansåg att Jörg Haider , som ordvrängare , har varit en röst för rasism och för främlingsfientlighet .
Han är en man som spelar på rädsla och som har utnyttjat människors sårbarhet .
Det är därför denna debatt är viktig - att markera att när man integrerar extremism händer något mycket omvälvande i Europa i dag .
( Applåder ) Jag skyndar mig att tillägga att vårt gräl inte gäller det österrikiska folket .
Vi respekterar det österrikiska folkets rätt till sin egen demokratiska process .
Vi försvarar det österrikiska folkets rättigheter och konstitutionella privilegier , men vi här i Europaparlamentet har en skyldighet att påminna oss om våra grundläggande principer enligt artikel 6 i fördraget - principerna om frihet , demokrati och respekt för mänskliga rättigheter .
Varje rättänkande person i denna kammare anser att dessa är universella och odelbara principer utan hänsyn till färg , klass eller tro .
Vi måste värna om och försvara dessa rättigheter och samtidigt tala om för det österrikiska folket : vårt gräl gäller inte er .
Beträffande det portugisiska ordförandeskapets initiativ vill jag framföra att vi stöder andemeningen och det politiska syftet bakom det .
Det är kanske inte ett perfekt initiativ i dess utformning men vi inser , herr ordförande , att dess grund är idealism och av det skälet är vi benägna att stödja det .
Jag delar ordförande Prodis uppfattning att gemenskapens metod är att föredra och vi måste titta på artiklarna 6 och 7 i fördraget .
I artikel 7 nämns möjligheten till tillfällig uteslutning i händelse av allvarliga och återkommande brott mot våra grundläggande principer .
Vi måste som institutioner hitta ett sätt att tillämpa och visa vad detta betyder , så att det får en verklig mening och innebörd .
Därefter kan vi arbeta tillsammans i enlighet med gemenskapens metod för att driva ut denna cancerböld mitt ibland oss .
Fru talman , jag vill säga några ord till Schüssel .
Schüssel är en man med ett hedersamt rykte i europeisk politik .
Han avser nu att rida in i regeringen på ryggen av en politisk tiger .
Herr Schüssel , ni tar på er ett mycket tungt , personligt , nationellt och europeiskt ansvar .
Det ansvaret , som ni herr Schüssel nu tar på er är att respektera ordalydelsen och andan i de europeiska fördragen .
Slutligen , fru talman , detta är en debatt som berör kärnan för våra demokratiska principer och institutioner och påminner oss om att priset för frihet är evig vaksamhet .
På denna kontinent , av alla platser , och mot bakgrund av vår erfarenhet av hatisk rasism som vi utstått tidigare och till så stor kostnad måste vi hävda att dagens debatt inte handlar om att hindra en stats suveräna rättigheter .
Det är ett hårdnackat krav från de demokratiskt valda i denna unions institutioner att vi som européer inte kan tillåta att man vrider tillbaka klockan .
( Livliga applåder ) Fru talman !
Det som händer i Österrike i dag är mycket allvarligt .
För första gången ställs Europeiska unionen inför risken att i ministerrådet , ibland oss , ha företrädare för ett parti som , uppenbarligen , uttalar sig och handlar i strid mot Europeiska unionens värderingar .
Jag vill göra tre kommentarer i frågan , för att illustrera problemets allvar .
Jag tror personligen att det handlar om ett första steg , om det nu äger rum , mot att banalisera extremisternas närvaro i regeringarna .
Jag tror också att det är en mycket negativ politisk signal till de sköra demokratierna i de länder som ansökt om medlemskap i Europeiska unionen .
( Applåder ) Jag tror slutligen att det är en politisk tillbakagång för Europeiska unionen som sådan , och därmed också en negativ signal utanför unionen , när vi talar i demokratins och de mänskliga rättigheternas namn .
Vissa har sagt att vi lägger oss i Österrikes inre angelägenheter .
Vissa har sagt att vi kritiserar det österrikiska folket och att vi faktiskt anklagar en framtida regering för ont uppsåt .
Är det att anklaga någon för ont uppsåt när man är uppmärksam på vad en politisk ledare säger sedan flera år och tydligt illustrerar en tendens som går tvärtemot allt det vi vill ?
Det är inte att anklaga någon för ont uppsåt och det är inte att kritisera det österrikiska folket när man talar vänligt till dem och säger : kära vänner , var uppmärksamma på vad som riskerar att hända hos er snart och sprida sig i hela Europa : inte någon brutal förändring - jag tror att Haider är alltför intelligent för det - utan en långsam erosion av de demokratiska rättigheterna , en långsam erosion genom kulturell spridning och detta är extremt farligt .
( Applåder ) Fru talman !
Tillåt mig att tacka er för ert inlägg i parlamentets namn .
Det var både relevant och politiskt intelligent .
( Applåder ) Jag skulle också vilja tacka rådets ordförandeskap för det strama , relevanta och behärskade inlägget .
( Applåder ) Och slutligen skulle jag vilja vända mig till det parti som , vare sig man vill det eller ej , är målet för våra uttalanden , nämligen PPE-DE .
Jag skulle vilja vända mig till Poettering och indirekt till Martens , som är en landsman och som varit vår kollega .
Herr Poettering !
Jag har hört att ni följer händelserna i Österrike .
Jag skulle ha önskat att ni föregrep dem och framför allt att ni i ert namns parti fördömde själva principen om en allians med människor som tillämpar verbalt våld , som kritiserar de svaga , håller främlingsfientliga tal och är tillmötesgående mot naziregimen .
( Applåder ) Herr Poettering !
Jag ifrågasätter inte er demokratiska oro , men jag tror att ni begår ett allvarligt politiskt misstag .
Och för att parafrasera en av mina ryktbara landsmän , Europas fader , Paul-Henri Spaak , skall jag säga att för er del är det inte för sent , men det är dags att ändra åsikt .
Fru talman !
I dag ställs Europeiska unionen enligt min grupp inför sin största politiska och etiska utmaning sedan den bildades .
Unionen har förvisso upplevt situationer där regeringen i ett medlemsland bestått av människor vars idéer och tillämpningar strider mot unionens värderingar .
Men med Haider och hans män är det den öppet rasistiska , antisemitiska och främlingsfientliga extremhögern som skulle vara med och besluta om vår gemenskap .
Att ingå i ett sådant framtidsperspektiv skulle , även om det sker under protest , innebära att man lovar att respektera en kraft som inte är respektabel .
Det skulle innebära att man banaliserar det oacceptabla i hela Europa , det skulle innebära att de högtidliga uttalandena från de europeiska institutionerna om de grundläggande värderingar som enar oss och som vi med rätta kräver att kandidatländerna skall respektera , förvandlas till värdelösa dokument .
Därför stöder vi andan i uttalandet från ordförandeskapet och fjorton medlemsländer , liksom det från Europaparlamentets talman då hon , till skillnad från kommissionens bleka och tvetydiga ståndpunkt , vill få oss medvetna om faran och åstadkomma en reaktion .
Det handlar naturligtvis inte för oss om att kasta skam över det österrikiska folket .
Alla åtgärder som vidtas skall ha den dubbla målsättningen för ögonen att förbjuda Haider utan att isolera det österrikiska samhället .
( Applåder ) Mer än någonsin behöver demokraterna i detta land vår solidaritet .
Den stora kraftsamlingen den 12 november förra året i Wien måste anpassas till den nya situationen .
Vi måste föra en dialog med dem , komma överens och verka vid deras sida , för att tillsammans bidra till att öppna ett annat perspektiv för det österrikiska folket.Slutligen måste vi också ställa oss frågan : hur har det kunnat bli så här ?
Det handlar förvisso för de österrikiska politikerna till att börja med om att besvara denna existentiella fråga för demokratins framtid , och börja med dem som nyss tagit den enorma risken att släppa fram extremhögern , men därutöver kan ingen , inbegripet Europeiska unionen , i våra ögon låta bli att ifrågasätta de anledningar som gör det möjligt för en skrupellös demagog att utnyttja den frustration och den rädsla som uppkommit genom en politik där alltför många befolkningar inte känner sig hemma .
Denna debatt ligger framför oss , men var och en av oss måste utan dröjsmål ta sitt ansvar .
( Applåder ) Fru talman !
Vi hade kunnat diskutera behovet av att stärka unionens grundläggande principer , för att kunna försvara dem gemensamt .
I stället är vi tvingade att debattera formella och reella fel som begåtts under dessa dagar .
Vi är chockerade över den politiska enfalden hos dem som med oförsiktiga ord har stärkt Haider i Österrike och förlöjligat unionen genom att trampa på fördragets artikel 7 och tillkännage okonstitutionella åtgärder .
Vi har aldrig någonsin varit vittne till en så allvarlig och klumpig inblandning i en medlemsstats interna angelägenheter .
Naturligtvis får man inte svika de idéer som ligger till grund för Europeiska unionen , och i det sammanhanget har den italienska regeringschefen förklarat att dessa principer står upptagna i ett fördrag : han nämnde Köpenhamnsfördraget , som jag - och alla ni andra - inte känner till eftersom det inte finns .
Kanske menade han Amsterdamfördraget , där ett antal principer räknas upp i artikel 6 och i artikel 7 anges förfarandet för att fastställa om en medlemsstat gjort sig skyldig till grava och upprepade kränkningar av de principer som anges i artikel 6 .
Men hittills förekommer inte någon kränkning , vare sig allvarlig eller upprepad , från Österrikes sida .
Förutom att vara en inblandning är ordförandeskapets uttalande diskriminerande , för den tillåter att man straffar ett folk och fråntar det rätten att välja vem man skall rösta på .
Hittills har vi inte sett någon politisk sammanhållning , inte ens i kampen mot den organiserade brottsligheten , eller för att försvara folkmordens offer .
Vi har inte skapat en gemensam valuta med ett minimum av stabilitet eller en ekonomi som gör att man verkligen lyckas bekämpa arbetslöshet och fattigdom .
Men på en enda minut har vi med en bildstormares ursinne lyckats förstöra unionens trovärdighet .
Sanktioner kan utdömas efter det att fördragen har kränkts och inte om ett demokratiskt valt parti bildar regering .
Hur skulle vi annars ställa oss till de kommunistiska stater där kommunisterna nu är på väg tillbaka : skall vi kasta ut dem också ur unionen om de kommer till makten , eller skall allt vara förlåtet för Stalins barnbarn ?
( Applåder från höger ) Det är med diplomati , övertalning , kultur , solidaritet , och inte med hot , som institutionerna kan få respekt och göra så att principerna respekteras , inte med antikonstitutionella medel .
Bilaterala förbindelser berör staterna , varför de 14 inte har med detta att göra .
Detta är att trampa på de europeiska institutionerna för att försvara politiska resonemang med en inkompetens som är värdig partier som just släppts fria ur totalitära system , men inte dem som företräder demokratiska traditioner .
Det är mycket , alltför mycket , som skiljer oss från Haider - vilket vi redan har skrivit flera gånger - bland annat hans anspråk på det italienska Alto Adige .
Men detta vet vi redan .
I dag får vi bittert lära oss att även andra företrädare för unionen inte längre stöder unionens demokratiska ansträngningar .
Vi är för legalitet och den demokrati som folken uttrycker , för respekt för den nationella suveräniteten , så länge den inte kränker fördragets principer eller de mänskliga rättigheterna .
Vi tror på Europa , medan andra verkar ha inlett arbetet med att montera ned unionen .
Detta är resultatet av en alltför snabb utvidgning och bristen på klarhet när det gäller roller och skyldigheter .
Vi har förverkligat ett Europa som bara utgörs av en skakig marknad , inte ett Europa av principer , av rättigheter och politik .
Och här ser vi konsekvenserna !
Allt vi kan göra är därför att uppmana kommissionen att fortsätta spela rollen av modererande kraft och ge uppmuntran åt dem som arbetar på att det österrikiska folkets självständighet och suveränitet skall få fortleva , så att det folket kan fortsätta att vara fritt och solidariskt gentemot andra folk .
( Applåder ) Fru talman , kära kolleger !
I dag är det hyckleriet som står på dagordningen .
Vi har ett råd som lyckats strunta i fördraget och använda en metod som helt ligger utanför artikel 6 och 7 och som , vid fall av allvarliga och långvariga brott , gör det möjligt att döma en stat .
I detta fall föreligger inte allvarliga och långvariga brott i Österrike .
Det finns risker - det är vi alla medvetna om - men det förekommer absolut för närvarande inget som helst vare sig allvarligt eller långvarigt brott .
Om man skulle tillämpa kriterierna i artikel 6 och 7 , om man skulle tillämpa kriterierna från Köpenhamn på våra institutioner , på Europeiska unionen , skulle denna europeiska union mycket sannolikt inte kunna bli medlem , på det sätt som man kräver av länderna i Central- och Östeuropa .
Och om vi talar om allvarliga och långvariga brott , kan vi kanske tala om vissa medlemsstater , vi kan tala om Italien och Frankrike , det första respektive tredje land som dömts av Europarådet , av domstolen i Strasbourg .
Vi kan , kära belgiska kolleger , tala om Belgien , om Dutroux-affären , tiotals och åter tiotals barn som rövats bort , torterats , våldtagits och mördats av personer från detta land och där undersökningarna fortfarande har kört fast .
Kära kolleger !
Vi skulle med en tredjedel av ledamöterna kunna tvinga rådet och kommissionen att ifrågasätta detta .
Vi skulle själva kunna ifrågasätta det faktum att österrikarna förkastar tio år , tretton år av " partikrati " som korrumperat och fått ett land - Österrike - att ruttna på samma sätt som det är på väg att korrumpera och låta länder som Italien , Belgien och andra av unionens medlemsländer ruttna .
Kära kolleger !
Vi skulle verkligen kunna fråga oss varför 76 procent av de belgiska medborgarna inte har något förtroende för rättvisan i sitt land , 56 procent av de franska medborgarna inte har något förtroende för rättvisan i sitt land och 53 procent av de italienska medborgarna absolut inte har något förtroende för sin rättvisa ...
( Talmannen avbryter talaren . )
Fru talman !
Min grupp , EDD , och i synnerhet mitt parti , är mycket oroade av denna debatt .
Vi kan inte stödja och vi stöder inte på något sätt Haiders åsikter och politik och vi beklagar hans hänvisningar till Tredje riket .
Men vi beklagar dock det faktum att ert parlament överväger att blanda sig i en vald regerings politik i något som helst land , särskilt ett som är en del av Europeiska unionen .
Mitt parti hemma är verkligen inte rasistiskt , men vi godkänner inte Europeiska unionens princip eller inblandning så lätt .
Kommer ni att blanda er i politiken i Storbritanniens parlament om vi blir valda ?
Fru talman !
Österrikes folk har talat genom att välja Haider till sitt parlament .
Jag tror de gav honom 28 procent av rösterna , så det kommer att bli en koalitionsregering .
Fru talman , får jag föreslå att ert parlament väntar och ser om Haiders parti kommer att påverka det landets politik .
Då och först då kan ni bedöma om mänskliga rättigheter påverkats .
Ert parlament kan överväga lämpliga åtgärder för att lösa den situationen och då , fru talman , först då kan ert parlament överväga att blanda sig i konstitutionella frågor i ett av Europeiska unionens länder .
Fru talman , som ledamot från det österrikiska liberala partiet respekterar jag den oro som vissa kolleger känner för den demokratiska utvecklingen i Österrike .
Ni kanske förvånas över min reaktion när jag säger att jag förstår att man är särskilt känslig och ifrågasätter Österrikes respekt för de mänskliga rättigheterna och dess ansvarskännande gentemot det egna förflutna och i fråga om den demokratiska stabiliteten i landet .
Österrike måste själv ta ansvaret för den ofta tvivelaktiga image som det med rätt eller orätt har i utlandet .
Våra regeringars vägran under många år att erkänna vår delaktighet i andra världskrigets fasor , och deras vägran att rättmätigt gottgöra de judiska offren och tvångsarbetarna , har väsentligt bidragit till denna negativa bild .
Nu har detta FPÖ ( Österrikiska liberala partiet ) på grund av det uppdrag de fick vid valet den 3 oktober 1999 , när den gamla regeringen valdes bort , gått in i en regeringskoalition med ÖVP ( Österrikiska folkpartiet ) .
Detta är den rättighet som medborgarna i en stat har , eftersom det är grundprincipen i en demokrati .
Efter att samtalen mellan SPÖ och ÖVP misslyckats försökte socialisterna bilda en minoritetsregering och bad FPÖ om deras stöd .
Vi erbjöds tre ministerposter - det kan ni se i tidningarna - just detta parti som här betecknas som fascistiskt !
När vi plötsligt avvisade detta erbjudande , började en våldsam hets och propaganda , som vi hittills inte kunnat förstå .
FPÖ är ett parti som länge varit etablerat inom den österrikiska politiken .
Det tillsätter ministerpresidenten i ett av de nio förbundsländerna och deltar i alla andra regeringar .
Varför , frågar sig många österrikare i dag , tolkas deras demokratiska beslut plötsligt som ett uttryck för en fascistisk inställning , varför har hetsen börjat just när de liberala avvisade stödet från en socialdemokratisk minoritetsregering ?
Här ägnar man sig åt ett fördömande som gör den hemskaste epoken i den europeiska historien till ett politiskt spektakel - utan att gå in på vårt program .
Det äcklar mig , när några av våra motståndare utnyttjar miljoner människors död i koncentrationslägrens gaskammare till billig propaganda , vilket exempelvis den italienske ledamoten Bertinotti gjorde , när han i går i italiensk TV anklagade Haider för att förneka förintelsen .
Ni borde skämmas , herr kollega !
Även om alla era politiska argument tar slut , har ni inte rätt att använda de mördade personerna för er billiga propaganda .
Ni förvandlas här inte till någon antifascist när ni betecknar en demokratiskt vald politiker som nazist !
Tvärtom , ni hånar de verkliga offren för nationalsocialismen och bagatelliserar de fascistiska diktaturerna .
Ni agerar på grund av era egna fördomar , ni avstår från all politisk diskussion och agerar just på det sätt som ni påstår att ni bekämpar .
Attacken mot Österrikes nya regering , försöket att påverka politiken i ett medlemsland är en förolämpning av den österrikiska befolkningen .
Därför är vi tacksamma för kommissionens speciella hållning .
I de nya koalitionsavtalen handlar det om en demokratireform , oppositionens rättigheter och plikten att lämna skadestånd åt tvångsarbetarna .
( Talmannen avbryter talaren . )
Fru talman , ärade kolleger !
Till att börja med vill jag fullständigt klarlägga en sak : Det finns i Österrike ingen risk för att det skall återuppstå något enpartisystem eller totalitärt system med högerinriktning .
Österrike är en stabil demokrati , där de mänskliga rättigheterna och friheterna garanteras av författningen och skyddas av ett oberoende rättsväsende .
Österrike är ett öppet land , där främlingsfientlighet och diskriminering inte hör hemma .
Det som pågår i Österrike är ett fullständigt normalt förfarande med en växling vid makten efter demokratiska val , där det gamla systemet valts bort och där man sökt och funnit en stabil parlamentarisk majoritet för de nödvändiga ekonomiska och sociala reformerna .
Det kommer att finnas en fungerande majoritet , liksom en fungerande opposition .
Det österrikiska folkpartiet , som jag företräder i detta parlament , var och är ett parti som alltid konsekvent har engagerat sig för att integrera mitt land i EU och som känner djup samhörighet med värdegemenskapen i Europeiska unionen , liksom med dess politiska principer för fördjupning och utvidgning .
Vi respekterar och accepterar diskussionen och kan också förstå den oro som uttalas i många av våra medlemsländer beträffande Österrikes framtida väg .
Vi har förståelse för det eftersom vi vet att vi på grund av vår historia för inte så länge sedan också har ett särskilt politiskt ansvar i samtiden .
Vårt land var inte bara det första offret för Hitlers diktatur , många var också gärningsmän , även om jag tillbakavisar all kollektiv skuld .
Österrike har , inte minst tack vare ÖVP , funnit sin väg in i Europeiska unionen .
Mitt land har sin plats inte utom utan inom Europeiska unionen .
( Applåder ) , och detta med alla rättigheter och skyldigheter !
Också en kommande regering måste därför bedömas efter vilka värderingar och principer den bekänner sig till i sitt regeringsprogram , och inte efter hur den fördöms , dels av politiska kontrahenter , dels av internationella medier .
Att bekänna sig till de mänskliga rättigheterna , demokratin och rättsprinciperna , till en uppriktig bearbetning av Österrikes roll i det förflutna , till vidarebefordran av information om mänsklighetens största brott under 1900-talet , förintelsen , kommer också att ingå i den grundläggande förståelsen hos en kommande koalitionsregering mellan ÖVP och FPÖ .
Mitt parti kommer att vara en garant för att mitt land bibehåller den Europapolitiska kursen och stannar kvar på den europeiska värdegemenskapens fasta mark !
( Applåder ) Fru talman , herr rådsordförande , ledamöter av kommissionen !
Detta är en svart dag för Österrike och för Europa .
Det kan inte heller Sichrovskys lögnaktiga konstruktion eller Stenzels lugnande ord ändra på .
Ty det har gått så långt att två oansvariga politiker , sönderslitna av maktsträvanden , säljer ut Österrikes image , dess politiska roll och delvis också dess ekonomiska intressen !
( Applåder , tillrop ) De byter ut detta mot en ställning som regeringschef och deltagandet i en regering .
Att Österrike förvandlas från ett aktat till ett utstött land finner de sig i , och även den isolering som hotar landet och därmed också delvis dess medborgare .
Jag anser - på samma sätt som många som i flera år kämpat mot Haider och hans politik , även mina kolleger i den socialdemokratiska delegationen här i kammaren - att alla åtgärder som vidtas av det internationella samfundet väger tungt och även är opassande , såvida de inte syftar på regeringen och dess företrädare .
Men min kritik - och det säger jag öppet - min vrede riktar sig uteslutande mot dem som har orsakat dessa reaktioner , herrarna Schüssel och Haider och deras partier , ( Applåder ) inklusive deras företrädare i detta parlament .
Kollega Poettering , detta är intressant : Ni befinner er i dag nästan i samma svåra position som jag , även om det är av andra anledningar , ty ni måste försvara något som ni inte vill försvara .
Ni försvarar en herr Schüssel - ni måste tänka på Schüssel i dag , som , efter vad jag hört , för kort tid sedan inte heller inbjöds till toppmötet med företrädarna för kristdemokratiska partiet .
Nu är argumentet , som även kollegan Poettering har använt , att Haiders förtrollande förmåga bara kan försvinna om han integreras i det politiska systemet .
Men jag påstår att han lika litet som andra högerextremistiska rörelser kan integreras i vårt politiska system och i detta Europa .
Den som livnär sig på fördomar mot utlänningar och minoriteter och som ger näring åt dessa fördomar , den som har inskränkthet och antiliberalism på sitt program , den som beter sig knölaktigt och arrogant i de internationella förbindelserna , och den som aldrig entydigt och otvetydigt har distanserat sig från nationalsocialismen , han är inte beredd att integreras och har inte för avsikt att bli det !
( Applåder ) Det är de konservativas stora historiska skuld att de frivilligt går till sängs med vargen och väntar tills de blir uppätna .
På så vis frodas vargen - även om ÖVP måste offra sig själva - i stället för att hållas stången .
Jag förstår att Europa och den civiliserade världen vill ha så litet som möjligt att göra med en sådan regering .
Men det finns också detta andra Österrike , detta Österrike som för x-tusende gången har demonstrerat mot att FPÖ skall delta i regeringen , och som kommer att fortsätta att demonstrera mot denna regering .
Jag ber detta Europa att stödja och hjälpa detta Österrike !
( Applåder ) Ju starkare detta Europa blir , och ju mer vaksamt det är mot auktoritära tendenser i Europa , desto mer framgångsrikt kan vi bekämpa högerextremismens rötter .
Ty Europa är och förblir den starkaste garantin mot främlingshat och demagogi eller rent av ett återfall i barbari .
Stöd det österrikiska folket mot denna regering !
( Applåder ) Fru talman !
Det här är ett historiskt ögonblick eftersom det nu äntligen står helt klart för oss alla att Europeiska unionen allt eftersom utvecklats till en värdegemenskap .
Vi inser detta nu när en medlemsstats regering håller på att få ett parti som veterligen inte respekterar dessa värden .
Jag vill också konstatera att de fjorton medlemsstaternas ställningstagande från rådets sida var berättigat , eftersom det här på sätt och vis också handlar om sammansättningen på Europeiska unionens regering , vilket gör att den här frågan angår även rådet .
Det är inte enbart Österrikes interna angelägenhet .
I egenskap av parlamentsledamöter måste vi särskilt betona att det arbete som inletts för att förstärka de grundläggande rättigheterna t.o.m. är viktigare än förut .
Det är viktigare än förut att respekten för och okränkbarheten hos de mänskliga rättigheterna samt minoriteternas rättigheter , alla de människors rättigheter som bor i Europeiska unionens område , är en väsentlig del av Europeiska unionens rättsstatsprincip , och därför måste också stadgan för de grundläggande rättigheterna göras juridiskt bindande .
Den får inte enbart förbli en förklaring .
Lika viktigt är det att stödja Österrikes demokratiska krafter , ingen av oss vill ju isolera Österrike .
Vi vet att majoriteten av österrikarna respekterar dessa värden .
De har också demonstrerat ; alla demonstrationer har inte ägt rum utanför Österrike .
Det är säkert också många väljare som röstat av protest , som länge velat ha en förändring i den österrikiska politiken .
Enligt min mening skall parlamentet stödja dessa demokratiska krafter .
Jag vädjar också till Österrikes president att han än en gång skall undersöka alla de möjligheter som finns att bilda en regering bestående av demokratiska krafter .
Fru talman , kära ledamöter !
Jag vill bara understryka värdet av den hållning som vår gruppordförande , Francis Wurtz , påminde om för ett tag sedan .
Jag uppskattar uttalandet från rådets ordförande och ståndpunkten från de 14 medlemsländerna som vägrar att ha officiella kontakter med den österrikiska regeringen så länge som Jörg Haiders parti ingår .
Det faktum att vi instämmer i detta blir desto viktigare eftersom vi , som bekant , har en kraftigt avvikande uppfattning när det gäller den politik som bedrivs av Europeiska unionen .
Detta gäller den ekonomiska och sociala politiken , det demokratiska underskottet , det faktum att unionens medlemsstater deltog i det dramatiska kriget på Balkan .
Detta vårt avståndstagande understryker ännu mer betydelsen av vårt instämmande i dag : det är något exceptionellt , för faran för att ett irrationellt och neonazistiskt parti återuppstår i Europa är exceptionell .
Den risken gäller inte bara Österrike , den gäller hela Europa .
Vi talar om oss själva , inte om Österrike .
Vi känner till de sociala faktorer som samverkar med arbetslösheten och osäkerheten , till att förstärka tendenserna i den riktningen .
Vi känner till de kulturella orsakerna - främlingsrädsla , rasism - men vi kan inte avstå från att i oförmågan och den bristande viljan från extremhögerns sida göra upp med nazismen och peka på risken för att det uppkommer en explosiv blandning i Europa .
Jag talar om Alperna , om alla våra länder .
Vi håller på att skapa förutsättningar som kan leda till att det uppkommer en fara för demokratin och det europeiska samhället .
Ordförandeskapets uttalande visade att man är medveten om det dramatiska i situationen .
Europa visar att man inte har glömt Auschwitz .
Europa möter ett spöke .
Men nu måste vi vara konsekventa i våra handlingar , och den första att vara konsekvent borde vara kommissionen , som i stället här har visat prov på en oklarhet och en brist på stadga som gör ordförandeskapets ståndpunkt ännu mer värdefullt .
Detta är den ändring vi måste kräva i kommissionens åtgärder .
Fru talman , kära kolleger !
I den grundläggande demokratiska principen om respekt för de mänskliga rättigheterna och folkens frihet och suveränitet , mot all gammal eller ny fascism , nazism eller kommunism , och med tanke på att samtliga föregående talare har talat om det österrikiska folkets suveränitet , så ser vi i dag hur denna suveränitet förnekas av just detta parlament .
När man läser det österrikiska liberala partiets partiprogram så finner man där ingenting som rättfärdigar anklagelserna om ett attentat mot principerna om frihet , demokrati och respekt för de mänskliga rättigheterna , de principer om grundläggande friheter och om rättsstaten som framhålls i artikel 6 i unionsfördraget .
Låt mig i stället rikta er uppmärksamhet på det faktum att den tjänstgörande ordföranden , som var så kritisk när det gäller Österrike , nyligen överlämnat invånarna i Macao till den demokratiska kinesiska folkrepublikens överhöghet .
Men kanske är det i dag , för att stärka demokratin inom unionen , lämpligt att isolera Österrike , kriminalisera ett parti som valts på demokratisk väg av det österrikiska folket och i stället släppa in det Turkiet som styrs av de grå vargarna i Europa .
Fru talman , ärade ledamöter !
Det är en högst allvarlig fråga vi diskuterar .
Det handlar om inte mindre än närvaron av en politisk makt i en medlemsstats regering , en makt vars lärosatser och principer är oförenliga med unionens föreställningar och moral som är heliga i de fördrag som unionen bygger på .
En genomläsning av artikel 1 i kapitel 4 i det österrikiska populistiska partiets program kan uppröra vilken demokrat som helst .
Accepterandet av den etniska gruppen som en avgörande faktor för en nation och påståendet att en folkgrupp är överlägsen alla andra , så som det påstås där , väcker gamla spöken till liv från ett århundrade som vi just har lämnat bakom oss , och som av vissa historiker betecknas som skräckens århundrade , en skräck som till vår bestörtning åter aktualiseras av den oacceptabla filosofin i Haiders politiska program .
Naturligtvis är det österrikiska folket ett självstyrande folk och naturligtvis skall vi respektera principen om icke inblandning i en medlemsstats inre angelägenheter .
Men det är inte det som är problemet .
Problemet är huruvida unionen kan förbli likgiltig inför bildandet av en regering i en medlemsstat , där ett parti med sådana drag ingår .
Vårt svar på denna avgörande fråga är nej .
( Applåder ) Bortom alla strategiska och taktiska överväganden , bortom alla eventuella rättfärdiganden som man gör på grund av främmande beteenden , bortom allt sådant , och oberoende av partiintressen och valtider , vill den spanska delegationen inom Europeiska folkpartiets grupp i parlamentet , helt i överensstämmelse med det spanska folkpartiet och Spaniens regering , uttrycka sitt stöd för uttalandet av rådets portugisiska ordförandeskap den 31 januari , vad beträffar dess innehåll , ton och konsekvenser .
( Applåder ) Konrad Adenauer sade vid något tillfälle - och han visste vad han talade om - att det säkraste sättet att lugna ned ett odjur är att låta dig slukas .
Historien är en provkarta på sådant som hade kunnat undvikas .
Därför , fru talman och kära kolleger , måste unionen och detta parlament ge tydliga signaler om att vi avvisar detta intoleransens , främlingsfientlighetens och totalitarismens odjur , för att bara nämna några av de misstag på den långa lista över avsägande av ideal , avståenden och opportunism som markerat Europas förflutna och som vi har fått betala ett högt pris för .
( Livliga applåder ) Fru talman , kära kolleger !
Vår union konstruerades kring tanken : " detta får aldrig hända igen " , och detta betydde " aldrig mer främlingsfientlighet , läger , antisemitism , aldrig mer någon bitter nationalism eller några krig " .
Europeiska unionen har inget annat syfte än viljan att överträffa denna fruktansvärda historia från det tjugonde århundradet som , i hjärtat av Europa , dödade hela idealet om humanism och som i dag fortfarande är högst aktuellt .
Det är inte sant när man säger att när en regering bildar allians med nyfascister , någonstans i Europa , är det bara ett problem med nationell suveränitet .
Vår union är inte någon sammansättning av stater-nationer som gör arrangemang sinsemellan för att förbättra sitt öde .
Det är en ödesgemenskap där alla demokrater tillsammans , när det viktiga ifrågasätts , när värderingar ifrågasätts , måste stå enade för att finna lösningar så att misstagen inte återupprepas .
Vi måste ta lärdom av det förflutna .
Under trettiotalet valdes Adolf Hitler demokratiskt , även om det var med minoritet , många tyckte att det inte var så farligt och , herr Poettering , i mitt land ansåg ett antal män och kvinnor till höger , men kanske också på annat håll : " hellre Hitler än Folkfronten " .
De föredrog sina lokalpatriotiska trätor framför det viktiga , och katastrofen var ett faktum .
Vi måste reagera snabbt , kraftigt och enat .
Herr Poettering !
Jag skulle ha velat höra er tala till den österrikiske presidenten eftersom vi vet att han i dag är mycket generad över denna smutsiga allians som ingåtts av en regering .
Vi måste alltså reagera snabbt och kraftigt .
Naturligtvis innehåller fördraget en spärr när handlingarna blir outhärdliga , och jag höll nästan på att säga " irreparabla " .
Historien har lärt oss att fascisterna börjar med att ge ros och ris : först ris , i de populistiska och främlingsfientliga talen , och sedan ros för att göra sig presentabla i institutionerna och successivt infiltrera dem , fördärva dem , ända till den dag de skrider till handling .
Och den dagen är det för sent .
Fördraget innehåller därför spärrar ; men vi är inte där ännu ; i dag måste vi förhindra att vi kommer så långt som till dessa spärrar .
Vi måste därför finna en politisk lösning .
I det stöder jag rådets förslag och jag beklagar en viss ömtålighet , en viss slapphet från kommissionen som ändå borde vara beslutsamt vaksam dag för dag , för fascisterna räknar med demokratins slapphet , de räknar med tiden för att slita ut oss och de hoppas slutligen kunna göra sig gällande .
Vi måste därför reagera snabbt .
Om vi i dag inte starkt stöder rådet kommer historien att döma oss och säga : de har genomfört ett politiskt München .
Fru talman !
Jag gläder mig över att den stora befolkningsmajoritetens vilja respekteras i Österrike och att , ur min synpunkt , demokratin vunnit en mycket viktig seger i och med den här regeringsbildningen .
Det måste stå alldeles klart : ett Europa som utvecklas som en sorts " Big brother " som på stalinistiskt sätt och med stalinistiska metoder vakar över vänsterns political correctness i den ena eller den andra medlemsstaten , ett sådant Europa undanber vi oss verkligen .
Den europeiska demokratin och den österrikiska demokratin behöver inte ta emot lektioner från någon annan och särskilt inte från en belgisk regering , till vilken av vapenhandlare finansierad korruption hör .
En belgisk regering som utsett ordföranden för ett sådant av domstolarna korruptionsdömt parti till ledamot av Europeiska kommissionen .
Vi tackar i dag Österrikes befolkning för den här demokratiska segern som är viktig för alla folk i Europa och för var och en som förespråkar frihet och yttrandefrihet .
Fru talman !
Denna debatt öppnades av Da Costa som bara bekräftar att EU : s ordförandeskap försöker påverka regeringssammansättningen i en medlemsstats regering .
Denna debatt och bakgrunden till den förstärkte åsikten att rådet , kommissionen och själva detta parlament domineras av socialister .
Min delegation som består av 37 konservativa och unionistmedlemmar från Förenade kungariket förkastar helt det österrikiska liberala partiets bakomliggandefilosofi , program och karaktär .
Vi delar den allmänna upprörelsen över dess inställning till historien , i synnerhet andra världskriget , men även dess politiska inställning till utvidgningen , invandring , rasfrågor och dess inställning till själva Europeiska unionen .
Men vi var också upprörda över vänsterns överseende med tyranniet , terrorn och övergreppen i f.d.
Sovjetunionen .
Även i dag är det verkligen hög tid för partiet av europeiska socialister att bryta de broderliga förbindelserna med Kinas kommunistparti .
Inte ett ord sades av dessa samma EU-regeringar om koalitionsregeringar med kommunistsympatisörer i franska eller italienska regeringar eller i regeringar i tyska stater eller till och med den brittiska regeringens beredvillighet att befordra personer med terroristanknytningar till ministrar i Nordirland i dag .
Detta , fru talman , är vänsterns skenhelighet .
Således fördömer vi den skenheligheten och dubbelmoralen , särskilt hos den brittiska regeringen och hos de andra huvudsakligen socialistiska ledarna i EU-regeringar och inkluderar även Förenta staternas .
Vi bör dock inse att den demokratiska processen ibland skapar obekväma resultat .
För detta krävs åtgärder för att ta itu med de bakomliggande orsakerna , däribland en granskning av själva valprocessen .
Det bör vara vår uppgift , inte politiskt ställningstagande .
( Applåder ) Fru talman , rådets företrädare , herr kommissionär !
För en vecka sedan avslutades i Stockholm den stora internationella Förintelsekonferensen .
Dess syfte var att bekämpa glömskan och det onda i dagens samhälle som uppträder i form av främlingsfientlighet och nynazism .
Det vore ett hån mot idén bakom denna konferens och hela det internationella samfundet att i dessa tider inbjuda ett nazistflirtande och främlingsfientligt parti i EU : s institutioner .
För det andra vill jag säga att vi måste vara konsekventa mot oss själva och våra värderingar .
Vi kräver av kandidatländerna och av samarbetsländerna i Loméavtalet att de skall respektera mänskliga rättigheter och visa tolerans gentemot nästan .
Vi måste göra detsamma mot oss själva .
Det är därför vi reagerar mot detta smusslande som pågår i Österrike .
Det går inte att fortsätta som om ingenting har hänt .
Vi står inför en vattendelare i unionen .
Unionen är inte bara en ekonomisk gemenskap , utan det är en värdegemenskap som vi tar på allvar .
Någonting har hänt : Unionen håller på att få ryggrad och själ .
Fru talman !
Alla har sagt det , det är en mycket viktig dag , det är dagen för den första debatten i det europeiska politiska livet .
Och det är ingen tillfällighet .
Det förefaller mig som om det möte vi har i dag inte är Europas möte , våra institutioners möte , med Österrike eller Haiders parti .
Det är Europas möte med sig självt , med dess existensberättigande , med anledningarna till att vi är närvarande här i kammaren .
Denna kammare finns inte till för varorna eller för pengarna .
Den och de europeiska institutionerna har byggts upp för värderingar , för moral och för en själ .
Men vi har under det tjugonde århundradet upplevt att demokratierna kunde hotas och att moralen , värderingarna och själen som jag nämnde kunde drabbas av ett dödligt virus som har ett namn : nationalistiskt förhärligande , populism och rasens överlägsenhet .
Och det räcker med att läsa programmet från Haiders parti , FPÖ , för att man i varje kapitel skall hitta nationalistiskt förhärligande , populism och rasens överlägsenhet .
Jag läser bara en mening som min vän Vidal-Quadras läst före mig " fosterlandet definieras genom sin plats , sin kultur och sin ras , såväl lokalt som etniskt och kulturellt " .
Vi kan inte acceptera sådana uttalanden .
( Applåder ) Om det finns någon mening med Europa och - jag ber om ursäkt att jag säger det till mina vänner - om det finns någon mening med den kristna demokratin , om det finns någon mening med den kristna demokratiska historien , måste den förklara sig radikalt oförenlig med påståendena i detta program och vägra , oavsett de utmärkta skäl som man framför varje gång som historien skickar runt fatet , att komma överens med denna typ av ideologi och denna typ av organisation .
Det är anledningen till att det förefaller mig som om Europaparlamentet , som är friare i sina handlingar och uttalanden än rådet eller kommissionen , måste välkomna dem bland staterna och de europeiska institutionerna som haft modet att säga " nej " , och som ni gjorde fru talman i vårt namn göra ett uttalande som ärar oss , och tydligt utan undanmanöver uttala sitt motstånd och sitt fördömande mot det som förbereds i Österrike , och att dagen för Münchenavtalet minnas uttalandet från en stor fransk demokrat som sade " när det handlar om att säga nej är det bästa tillfället det första " .
( Applåder ) Fru talman !
Vi är bekymrade .
Vi , det är de belgiska kristdemokraterna och lyckligtvis väldigt många andra kolleger med oss .
Den koalition som håller på att bildas i en av medlemsstaterna är absolut en österrikisk angelägenhet men det hela har utan tvivel även en europeisk dimension .
Vad binder oss samman i Europa .
I första hand värdena och principerna om frihet , demokrati och respekt för de mänskliga rättigheterna .
Ordföranden för det österrikiska liberala partiet , Haider , har flera gånger visat att han inte tillräckligt högt värderar ens de grundläggande formerna av diplomatisk artighet .
Han är en farlig man .
De kristdemokratiska partierna i mitt land har för länge sedan valt , och håller fast vid , att visserligen lyssna till de högerextremistiska väljarnas protester men att aldrig förhandla med de högerextremistiska ledarna .
Värden måste komma före makt .
Därför beklagar vi det som sker i Österrike .
Vi är till och med skakade av det .
Vi är mycket besvikna .
Vi uppmanar ÖVP att i sista hand ändå undersöka andra lösningar .
Vi fortsätter att påminna om artikel 6 i fördraget .
Vi fortsätter kämpa mot banaliseringen av den extrema högern .
Om koalitionen ändå blir av så uppmanar vi våra kolleger i ÖVP att både i program och i ord och handling garantera att de principer och värden som utgör grunden för den europeiska integrationen respekteras .
Fru talman , mina damer och herrar , kolleger !
Det vilar ett stort ansvar på Österrike .
Fru talman , mina damer och herrar !
Det är uppenbart att vi i detta parlament i stor utsträckning är överens när det gäller att avvisa Haider och hans politik , men det är också klart att vi har olika uppfattning om hur man på effektivaste sätt skall kunna bekämpa denna politik .
Har ni tänkt på vad debatten här och uttalandet från rådets ordförandeskap förra veckoslutet får för effekt i Österrike ?
Har ni någon gång frågat er om vi inte också är ansvariga för den fortsatta utvecklingen av det politiska läget i Österrike , om vi här sätter oss till doms över detta ?
Har ni någon gång frågat er vad som skulle ske om önskemålet från en kollega uppfylldes och val ägde rum i Österrike inom de närmaste dagarna ?
Enligt samstämmiga uppgifter från alla observatörer skulle Haider bli ännu starkare .
Vem kan vilja något sådant ?
Är det inte vårt ansvar att tänka över hur vi skall bekämpa denna politik ?
Europa är en rättsgemenskap .
Till de principer som vi skall företräda hör demokrati , aktning för de mänskliga rättigheterna och rättsprinciperna .
Till kravet om demokrati hör att man inte ogillar valresultat , utan måste respektera dem , och därför måste vi respektera om österrikarna , av orsaker som har med deras politik att göra , beslutar så som de nu har gjort .
Det är en rättsprincipiell fråga att rådets ordförandeskap inte får yttra sig så som det har gjort , på ett sätt som motsäger fördraget .
( Applåder ) Det är politiskt klokt att inte isolera ÖVP , utan stödja ÖVP som ett tveklöst demokratiskt , rättsstatligt och uppenbart europeiskt parti , så att Österrike lika tveklöst förblir en medlem av denna europeiska gemenskap , och därför måste ÖVP-kollegerna få vårt stöd i denna svåra situation , och isolering är absolut fel väg !
( Applåder ) .
( EN ) Fru talman !
Där jag kommer från säger man " en walesare har tre tillfällen " och tre gånger , vilket jag tror ni kommer att upptäcka under den debatten , framförde jag min önskan att kortfattat lämna synpunkt på vad som har varit en utmärkt och vid flera tillfällen känslig debatt .
Först och främst vill jag framföra mitt tack på ordförande Prodis vägnar och mina kollegors i kommissionen för det stöd och samförstånd som flera ledamöter av kammaren visade för kommissionens ståndpunkt i det uttalande som vi gjorde i går .
Jag måste naturligtvis även reagera på det faktum att man under debatten gjorde anspelningar på - och jag använder några av de ord som användes - tvetydigheten , eftergivenheten och vekheten i kommissionens yttrande .
Jag känner mig förpliktad att till denna kammare framföra att det finns ingen tvetydighet eller vekhet eller eftergivenhet i det yttrande som gjordes eller de åtgärder som kommissionen vidtog i denna fråga .
Vi hänvisade i vårt uttalande i går morse , liksom ordföranden gjorde i eftermiddags , uttryckligen till det faktum att vi delar den oro som fjorton medlemsstater framförde i sitt uttalande i måndags .
För det andra , påpekade vi i mycket specifika termer att vi kommer att arbeta nära och tillsammans med alla medlemsstater för att granska situationen och dess utveckling i Österrike .
För det tredje , vi förklarade mycket klart att vi utan rädsla opartiskt kommer att hålla fast vid principerna och bestämmelserna i artikel 6 i fördraget och att vi skall göra vad som ankommer på oss enligt artikel 7 i fördraget för att säkerställa att dessa principer för frihet och demokrati och grundläggande fri- och rättigheter upprätthålls .
Det finns alls ingen eftergivenhet , vekhet eller tvetydighet i något av detta .
Och när jag säger att kommissionen intog denna ståndpunkt innefattar jag min kära kollega Franz Fischler , som kommer från Österrike och som återigen bevisade sin integritet och sin oberoende ställning som ledamot av Europeiska kommissionen under ed genom att delta i det uttalande som vi gjorde i går morse .
Var och en som därför bjuder in Franz Fischler till sitt hem för att av någon anledning förklara det faktum att han är av österrikisk nationalitet bör granska sina egna motiv i samband med en debatt som nödvändigtvis har skymts av hänvisningar till främlingsfientlighet och även mer farlig ondska i denna värld .
Jag säger det i vänskap och vördnad för min vän och kollega Franz Fischler .
Får jag också tillägga , fru talman , att förståelsen hos ordförandeskapet , det portugisiska ordförandeskapet , för vår ståndpunkt mycket klart bekräftades av Da Costa när han sade , och jag citerar honom , att " Portugal och övriga medlemsstater önskar säkerställa att gemenskapsmaskinens arbete inte störs av den nuvarande situationen " .
Det är förvisso i allas intresse .
För att kunna garantera att fördraget efterlevs och att vi håller vad som beskrevs som gemenskapsmaskinen i gång följer vi det tillvägagångssätt som lades fast i vårt uttalande i går .
Vi skall fortsätta att göra det , fru talman , på ett opartiskt sätt .
Det är vår plikt .
Det är också en fråga om övertygelse .
Min sista punkt är följande .
Vi inser innebörden i denna viktiga debatt .
Det finns flera personer här som liksom jag själv under många år tidigare blivit vana vid Haiders stötande uttalande , främlingsfientligheten i många delar av hans politik och den strategi han utvecklat att omväxlande göra aggressiva uttalanden och sedan framföra ursäkter , ibland påföljande dag .
Vi inser det och vi kommer även ihåg det dåliga och selektiva minne han ibland visar om nazismen .
Och när vi minns det , som så många andra runt om i denna kammare , väcks naturligtvis mina och mina kollegors instinktiva känslor till liv .
Men kommissionen måste agera på grundval av värderingar och lagar och inte bara på grundval av instinkter .
Det är därför vi kom fram till vår slutsats i går morse .
Det är därför vi håller fast vi den slutsatsen medan vi fortsätter att upprätthålla principerna och lagarna .
Utan vekhet , utan eftergivenhet , utan tvetydighet men till nytta för hela unionen och varje medlemsstat i unionen och dess folk .
Vi skall fortsätta att göra det energiskt och konsekvent och som Cox sade i debatten , " ovillkorligen med hög bevakning " .
Jag undrar , då Da Costa har lyssnat till dessa inlägg långt bak i kammaren , om herr Kinnock kan bekräfta att kommissionen stöder den åsikt som Da Costa klart fastslog i dag och som även fastslogs i ordförandeskapets nyligen gjorda uttalande å regeringschefernas vägnar .
Stöder kommissionen rådet ? .
( EN ) Fru talman !
När kommissionen i går morse sade att den konstaterar att de åsikter som framförts vara ett gemensamt uttalande av fjorton medlemsstater och att den delar den oro som låg till grund för den åsikten , anser jag att det kan förutsättas att den sedan i går morse och så snart som kommissionen kunde diskutera frågan den haft samma åsikt som de fjorton medlemsstaterna .
Tack , kommissionär Kinnock .
Jag tror att vi upplevt en stor politisk debatt , i nivå med situationen och vad man kunde vänta sig .
Tack , kära kolleger .
Jag förklarar den aktuella och brådskande debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.00 .
 
Tillämpning av försiktighetsprincipen Nästa punkt på föredragningslistan är meddelande från kommissionen om tillämpning av försiktighetsprincipen . .
( EN ) Jag vill börja med att säga att jag är glad att få lägga fram detta meddelande om tillämpning av försiktighetsprincipen , och det har författats tillsammans med David Byrne och Erkki Liikanen .
Försiktighetsprincipen är inte ett nytt koncept .
Den har tillämpats av gemenskapen ganska länge nu på en rad politikområden som miljö , folkhälsa , djur- och växtskydd och den nämns uttryckligen i miljöbestämmelserna i EG-fördraget efter Maastricht .
Den återfinns även i en rad internationella texter , till exempel Rioförklaringen och allra senast i biosäkerhetsprotokollet .
Innebörden i försiktighetsprincipen är uppenbar .
Den handlar om att vidta åtgärder på ett bestämt politikområde när den vetenskapliga delen inte är klarlagd , men där det finns skälig grund till oro för att de potentiella riskerna är tillräckligt stora för att kräva åtgärder .
Tillämpningen av försiktighetsprincipen har emellertid fått en ökad uppmärksamhet under senare år .
Händelser som BSE och dioxinkrisen har stimulerat till en växande offentlig debatt om vid vilka omständigheter försiktighetsåtgärder är berättigade och nödvändiga .
Med hänsyn till detta ökande intresse ansåg därför kommissionen att det skulle vara lämpligt att lägga fram ett meddelande för att fastslå kommissionens ståndpunkt om användningen av försiktighetsprincipen .
Det finns två huvudsyften med meddelandet .
Dels att förklara på ett tydligt och konsekvent sätt hur kommissionen tillämpar och avser att tillämpa försiktighetsprincipen i sin riskbedömning , dels att fastställa riktlinjer för dess tillämpning baserade på motiverade och konsekventa principer .
Vi hoppas också att meddelandet skall bidra till att skapa en bättre allmän förståelse för hur risker skall hanteras och att skingra farhågor om att försiktighetsprincipen skulle kunna användas på ett godtyckligt sätt eller som en förvrängd form för skyddstullar .
Kommissionens utgångspunkt för att tillämpa försiktighetsprincipen är behovet att garantera en hög skyddsnivå på områdena , miljö , folkhälsa , djur- och växtskydd .
Naturligtvis kan denna målsättning inte användas för att rättfärdiga irrationella eller godtyckliga åtgärder , men det innebär att åtgärder fortfarande kan vidtas även i situationer där vetenskapen är oklar .
Medan försiktighetsprincipen inte innebär att man gör politik av vetenskap , vilket några har velat göra gällande , för den oss fram till vägskälet mellan vetenskap och politik .
Det inledande beslutet att tillämpa försiktighetsprincipen beror till stor del på den skyddsnivå som eftersträvas och den risknivå som beslutsfattare är beredda att godta för samhället .
Den är därför politisk till sin natur .
De åtgärder som senare kan vidtas måste självklart följa de allmänna principer som tillämpas för hantering av risker och riktlinjerna för att tillämpa försiktighetsprincipen är därför den viktigaste delen i dokumentet .
De åtgärder som vidtas skall stå i proportion till den valda skyddsnivån - det vill säga , vi använder inte en hammare för att knäcka en nöt .
De måste vara icke-diskriminerande i sin tillämpning , det vill säga , åtgärder bör inte skilja sig på grundval av geografiskt ursprung .
Och de måste överensstämma med redan vidtagna åtgärder .
Exempelvis om en produkt har blivit godkänd , bör likartade produkter också godkännas .
Åtgärder baseras på en granskning av eventuella fördelar och kostnader för åtgärder eller brist på åtgärd ; det vill säga åtgärderna skall vara kostnadseffektiva och kunna utvärderas mot bakgrund av ny vetenskaplig information och klart fastslå vem som är ansvarig för att lägga fram de vetenskapliga bevis som krävs för en mer djupgående riskbedömning , det är bevisbördan .
Alla dessa element skall tillämpas kumulativt .
Det är också viktigt att komma ihåg att det finns ett brett urval av åtgärder som kan vidtas vid tillämpning av försiktighetsprincipen .
Till exempel ett forskningsprogram , allmänna informationskampanjer , rekommendationer och så vidare .
Att tillämpa försiktighetsprincipen medför därför inte automatiskt ett förbud .
Det första meddelandet är inte avsett att bli det slutgiltiga ordet i denna fråga .
Men det är första gången som kommissionen har lagt fram ett strukturerat dokument om principen och dess tillämpning .
Genom att fastlägga någorlunda detaljerat hur kommissionen tillämpar och avser att tillämpa försiktighetsprincipen hoppas vi kunna klargöra situationen på gemenskapsnivå och att medverka i den pågående debatten på europeisk och internationell nivå .
Herr talman , fru kommissionär !
Tack så mycket för förklaringen .
Jag har tre mycket korta frågor .
Den första frågan : Vi har fått vänta mycket länge på ett enhälligt yttrande från kommissionen om försiktighetsprincipen , och tidigare har det över huvud taget inte stått klart om kommissionen talar med en röst .
Är det som ni i dag här har lagt fram också den åsikt som era kolleger med ansvar för industri , utrikeshandel , konkurrens och den inre marknaden har ?
Ni kommer säkert att säga ja , men jag vill få veta följande av er : Känner dessa herrar till vilka konsekvenser det får ?
Nästa fråga , fru Wallström : När kommer ni att börja att tillämpa detta i lagstiftningen , när det gäller exempelvis kemikalier eller lagstiftning på andra områden ?
Den sista frågan : Kommer vi att kunna urskilja var detta tillämpats i lagstiftningen ?
Det betyder : kommer det att finnas en extra sida i varje förslag som talar om att försiktighetsprincipen har tillämpats och att man kommit fram till detta resultat ? .
( EN ) Tack så mycket , Dagmar Roth-Behrendt , för dessa frågor .
Naturligtvis delas detta av hela kommissionen .
Detta är ett allmänt meddelande som skrevs av oss tre , David Byrne , Erkki Liikanen och jag själv , men det har godkänts enhälligt i kommissionen i dag .
Det fick starkt stöd från övriga kommissionärer och samråd om det har hållits i hela kommissionen .
Så vi har verkligen genomarbetat detta dokument och jag är säker på att de alla kan beskriva de riktlinjer och principer som fastslås i detta dokument .
Ja , jag kan säga att vi redan använder detta sätt att arbeta med olika , svåra frågor som en ny kemisk strategi till exempel .
Jag är också säker på att vi uttryckligen kommer att nämna den när vi arbetar med denna princip .
Vi har nyligen haft ett fall där vi använde försiktighetsprincipen när vi måste förbjuda phtalater i mjuka PVC-leksaker och naturligtvis använder vi den på flera olika miljöområden .
Den har framför allt använts på miljöområdet , men naturligtvis också när det gäller folkhälsan .
Så vi skall försöka vara mycket tydliga om hur och när den skall användas .
Herr talman , fru kommissionär !
När det gäller förhållandet mellan vetenskapen å den ena sidan och försiktighetsprincipen å den andra sägs det i meddelandet att det alltid krävs ett politiskt beslut för att använda försiktighetsprincipen när de vetenskapliga bevisen är bristfälliga .
På det sättet lägger man naturligtvis över en hel del makt i händerna på vetenskapen .
Man kan undra vilken sorts vetenskapsmän som kommer att lämna den dokumentationen och vad står de för ?
I meddelandet står också att om det finns en tillräckligt stor erkänd minoritet av vetenskapsmän så räcker det för att kunna hänvisa till försiktighetsprincipen .
Jag skulle vilja fråga , vad är då definitionen för en erkänd minoritet ?
Hur beskriver ni en sådan ?
Hur kommer ni fram till en erkänd minoritet ?
När det gäller det politiska beslutet så skulle jag också vilja fråga : vem fattar det politiska beslutet ?
Är det kommissionen ?
Är det rådet ?
I vilken utsträckning kommer parlamentet att kunna delta i det beslutsfattandet ?
Vilken funktion har den vetenskapliga kommittén ?
Vilken roll kommer inom kort den myndighet för livsmedel som ni skall inrätta att spela ?
Avslutningsvis , kommer hela beslutsfattandet att ske på ett öppet och genomblickbart sätt ?
Det är mina tre frågor . .
( EN ) Ja , herr talman , det är sant .
Det fanns många och svåra frågor och inte alltid kristallklara men jag skall försöka besvara några frågor .
Vem vill fatta beslutet , vilka är beslutsfattarna ?
Jo , det beror på vilka lagstiftarna är .
Detta är en del av riskhantering .
De måste granska exempelvis omsorg om människor i förhållande till en särskild fråga och de måste göra en bedömning mot bakgrund av vad som är känt om vetenskapliga bevis i ett bestämt fall .
Men det är sant att det krävs inte uppbackning av en stor majoritet av det vetenskapliga samfundet för att kunna använda försiktighetsprincipen .
Den kan tillämpas på basis av bevis från en minoritet eller när vetenskapliga bevis är ofullständiga .
Det är naturligtvis där som ni gör en avvägning mellan denna princip som ett politiskt verktyg och vetenskap .
Det är inte alltid lätt att beskriva exakt hur denna process fungerar , men det är inte tal om att förändra den vetenskapliga grunden .
Vi använder experterna för att få så mycket vetenskaplig information och fakta som möjligt innan vi fattar ett beslut - och det bör också ske i framtiden .
Ni måste betrakta denna princip som ett verktyg för riskhantering .
Ni måste besluta om ni vill utsätta människor för fara till exempel , eller om ni vill skydda miljön , och ni måste utvärdera de vetenskapliga bevis som finns tillgängliga .
Ni måste bedöma allt detta och utvärdera vad vetenskapen visar .
Därefter beslutar ni om att vidta en åtgärd eller inte , att göra något eller inte .
Således finns det inga svar på alla era frågor , men det förändrar inte det system med forskare som vi använder i dag , eller det system med experter som vi använder i dag .
Herr talman !
Jag har en fråga som gäller ett konkret och aktuellt fall , i vilket försiktighetsprincipen skulle kunna tillämpas .
Det gäller bromerade flamskyddsmedel .
Det är så att dessa ämnen nu upptäcks ; det finns ökade koncentrationer av dem i både människor och miljö .
Det finns många som hävdar att de medför stora risker , medan andra ifrågasätter hur stora riskerna är med dessa ämnen .
Nyligen uppmanade både Sverige och Danmark i ministerrådet kommissionen att ta ett initiativ för ett förbud mot bromerade flamskyddsmedel .
Jag undrar då om ni förbereder ett sådant förbud och om det inte skulle passa väldigt väl in i er syn på själva försiktighetsprincipen att komma med ett sådant initiativ . .
Herr talman !
Tack så mycket , Jonas Sjöstedt , för denna fråga .
Frågan om bromerade flamskyddsmedel är viktig .
Den väcktes alldeles nyligen i miljörådet av ett antal ministrar som vill att kommissionen skall titta på vad det finns för underlag och vad som kan behöva göras .
Vi är i färd med att se på denna fråga och bedöma vilka kunskaper vi har i dag och vad som är möjligt att göra .
Låt mig dock få påminna om att användning av försiktighetsprincipen inte behöver vara samstämmigt med att det skall bli ett förbud , ett totalförbud .
Det kan finnas en rad olika åtgärder som kan vidtas .
Därför skall det inte omedelbart tolkas som ett förbud .
Vad gäller de bromerade flamskyddsmedlen kan det så småningom ändå bli det , men det är viktigt att säga att försiktighetsprincipen tillåter att man använder hela spektrumet av politiska insatser och åtgärder .
Denna fråga är aktuell i allra högsta grad .
Kommissionen skall göra sitt jobb och titta ordentligt på den innan vi återkommer med en bedömning av vad som behöver göras .
Ni framförde att försiktighetsprincipen inte bör användas som ett förtäckt handelshinder .
Är denna uppfattning överensstämmande på båda sidor om Atlanten ?
Jag tror att vi kommer att få problem med i synnerhet hormonbehandlat kött och genetiskt modifierade grödor .
Kommer amerikanerna att ha samma uppfattning i denna fråga som vi ? .
Herr talman !
Jag är glad att kunna meddela att vi i Montreal precis har skrivit under ett protokoll om biosäkerhet .
Där lyckades vi enas i ett internationellt forum om definitionen av försiktighetsprincipen .
Jag anser att det är ett genombrott , att vi lyckades avsluta detta protokoll .
Jag tror att det kommer att bilda skola för framtida diskussioner om försiktighetsprincipen .
Vi kommer att kunna använda detta som ett exempel på hur man skall tolka försiktighetsprincipen .
Den är dessutom även accepterad som ett viktigt och verkningsfullt instrument .
Herr talman !
Jag har två frågor ; jag skall försöka fatta mig väldigt kort .
Den första frågan gäller genomförandet av försiktighetsprincipen .
Som jag har förstått det , har det varit vissa oklarheter om hur man skall uppfatta detta .
Är det så att man först skall göra en riskbedömning där man inkluderar en kostnads- och nyttoanalys , alltså en cost-benefit-analys ?
I så fall blir jag ganska orolig , eftersom det väl var meningen att man inte skall använda en cost-benefit-analys som ett redskap för att avgöra om man skall introducera försiktighetsprincipen , utan försiktighetsprincipen skall komma först .
Min andra fråga gäller bevisbördan .
Jag minns när Margot Wallström introducerades som kommissionär i utskottet .
Då var hon inne på att man skulle vilja ha en omvänd bevisbörda .
Det vill säga att tillverkaren av en produkt skall visa om den är farlig eller inte .
Jag vill veta om detta också gäller i det dokument som kommissionen har presenterat nu . .
Tack så mycket , Inger Schörling .
Detta är två viktiga frågor .
Det är bra att jag får tillfälle att klargöra dem .
Nej , man måste inte börja med att göra en cost-benefit-analys , utan detta skall baseras på en bedömning av vad vi vet , vad vetenskapen kan berätta för oss och hur vi skall se på det jämfört med de risker som vi bedömer finns för miljön eller för hälsan hos människor och djur .
Däremot när man har bestämt sig för att vidta en viss åtgärd , då bör man välja en kostnadseffektiv åtgärd , så att man faktiskt inte tar till åtgärder som är helt orimliga när det gäller effektivitet .
Det är alltså inte så att man måste börja med en cost-benefit-analys .
Den andra frågan rör den omvända bevisbördan .
Det är alldeles riktigt att vi behöver tillämpa det i vissa fall .
Jag har använt exemplet kemikaliestrategin som ett bra exempel på ett område där vi behöver göra detta .
Då handlar det emellertid om det sakområdet , medan man kan säga att detta meddelande om försiktighetsprincipen är horisontellt ; det gäller alla olika specifika politiska sakområden .
Därför diskuteras inte speciellt i detta sammanhang en omvänd bevisbörda eller hur bevisbördan skall se ut , utan det handlar i stället om det politiska beslutsfattandet och grunderna för detta .
Det är dock alldeles riktigt att vi t.ex. när det gäller kemikalier måste se till att vi får en omvänd bevisbörda .
Herr talman !
Jag anser att försiktighetsprincipen för att fungera måste tillämpas ganska radikalt , för annars förlorar vi oss i tolkningarnas irrgångar .
Låt mig ge ett exempel : det visar sig att en antikryptogam gör så att det föds blinda barn , medlet är med andra ord teratogent .
OK , detta är en antikryptogam , ett antimögelmedel .
Den teratogena effekten har påvisats av ett enda engelskt laboratorium , kanske det enda laboratorium som har gjort några undersökningar .
Jag anser då att försiktighetsprincipen , med tanke på att det rör sig om ett så allvarligt hot mot hälsan , kräver att produkten omedelbart skall förbjudas , så som till exempel Nya Zeeland har gjort .
Låt mig alltså ställa den här frågan : när människors hälsa står på spel , eller man riskerar allvarliga hälsoeffekter , skall man då kanske göra en kostnads / intäktsanalys ?
Den kostnad som ett blint barn innebär är enligt mitt förmenande alltför hög , det finns inga vinster som kan uppväga den .
Jag vill därför veta om försiktighetsprincipen i det här fallet , så som ni tolkar den , fru kommissionär , förutsätter att produkten under alla omständigheter skall tas ur marknaden till dess att bevis om motsatsen har framlagts av andra laboratorier . .
Herr talman !
Jag är den första att önska att vi kan tillämpa försiktighetsprincipen på ett sådant sätt att det upplevs som radikalt till skydd för människors hälsa och för miljön .
Det är klart att jag inte kan ta ställning till det speciella fall och den speciella produkt som nämns här , men jag skall direkt gå tillbaka och se vilken information jag kan få fram om just detta fall .
Sanningen är ju att väldigt många medlemsstater , förvisso också andra nationer , har vidtagit åtgärder för att skydda sin befolknings hälsa på ett sådant sätt att man har använt försiktighetsprincipen , även om man inte alltid har kallat det så .
Det är naturligtvis så att det inte i första hand är frågan om en kostnad ; det kan nämligen bli en enorm kostnad för samhället om man undviker att vidta en viss åtgärd .
Det får inte heller vara så att man sitter och räknar vad ett människoliv kostar gentemot att vidta en åtgärd .
Jag tycker dock att det är alldeles självklart att när det så småningom är dags att besluta sig för en åtgärd , är det ofta så att man har många olika handlingsalternativ .
Då skall man titta på vad som ger bäst resultat .
Jag kan inte låta bli att berätta om ett tillfälle när detta uttryck användes av personer som man kanske inte alls skulle kunna tänka sig använda ordet kostnadseffektiv , nämligen vid ett besök i Afrika .
På ett hospice för aidspatienter träffade jag två irländska , katolska nunnor som skötte om döende aidspatienter .
De var de första att säga att vi måste varje dag tänka på att göra det som är mest kostnadseffektivt , därför att det måste räcka till våra stackars patienter här ; vi måste vara mycket noga med hur vi använder resurserna .
Jag menar att vi kan lära oss något av detta .
Vi måste ju alltid se till att vi använder våra resurser på effektivaste sätt och så att de kommer till hjälp på bredast möjliga sätt .
Det är alltså inte korrekt att man först måste börja med någon sorts cost-benefit-analys , vilket också förklaras i detta meddelande .
Man skall titta på vad vetenskapen erbjuder för kunskaper , och man skall använda detta som ett viktigt politiskt instrument för att skydda miljön och människors hälsa .
Herr talman !
Det är en sällsynt nåd att få en andra möjlighet att ställa en fråga !
Fru kommissionär , jag vill än en gång komma tillbaka till min första fråga , som kanske lät skämtsam , när jag frågade efter de andra kommissionärerna .
Ni besvarade den också så som jag visste att ni skulle göra .
Jag skulle vilja knyta samman den med något som Goodwill frågade , nämligen med vårt förhållande mellan försiktighetsprincipen och världen utanför Europeiska unionen .
Jag frågar ju inte detta utan orsak .
Ni har med all rätt sagt att försiktighetsprincipen är nödvändig just när vetenskapen ännu inte har några bevis .
Hur skall vi se till att vi inte alltid blir möjliga att angripa , t.ex. av våra partner i USA - och då räcker inte bio safety-protokollet till ?
Hur skall vi se till att inte industripolitikerna och utrikeshandelspolitikerna sparkar undan benen för er på samma sätt som de tidigare alltid gjorde med era företrädare ?
Det är just det som det handlar om , annars behöver vi här inte tala om försiktighetsprincipen , fru kommissionär ! .
Herr talman !
Jag tycker att det är väldigt viktigt att visa på de riktlinjer som finns för användande av försiktighetsprincipen i detta meddelande som ett sätt att tillbakavisa påståendena om att vi alltid vill använda detta av protektionistiska anledningar .
Jag är säker på att vi kommer att få fler konflikter med t.ex.
USA .
Vi skall inte vara naiva och tro något annat .
Ända sedan vi skrev under detta protokoll i Montreal , har vi emellertid ett internationellt erkännande och en gemensam definition inskriven i ett protokoll som handlar om miljö , hälsa och handel .
Det utgör därför ett gott exempel .
Vi skall inte tro något annat än att det kan dyka upp konflikter även i fortsättningen , men nu kan vi visa att vi inte använder försiktighetsprincipen godtyckligt .
Vi har nu ett antal riktlinjer för detta , och vi har ett starkt stöd hos våra respektive befolkningar för att använda försiktighetsprincipen , vilket tydligt fastläggs i detta meddelande .
Tack , fru kommissionär .
Den uppmärksamhet som ägnats åt den politiska försiktighetsprinipen har lett till att vi har diskuterat frågan i ungefär två timmar och nu anses den frågan så att säga ligga utanför den normala rutinen , även om , som vi har kunnat konstatera av de inlägg vi har hört i dag , från frågorna och svaren , det är en fråga som man fäster stor vikt vid .
Jag förklarar debatten avslutad .
 
Regeringskonferensen Nästa punkt på föredragningslistan är betänkande ( A5-0018 / 2000 ) av Dimitrakopoulos och Leinen för utskottet för konstitutionella frågor om sammankallandet av regeringskonferensen ( 14094 / 1999 - C5-0341 / 1999 - 1999 / 0825 ( CNS ) ) . .
( EL ) Herr talman !
Jag skall till att börja med tacka det portugisiska ordförandeskapet och kommissionen för alla de mycket nyttiga kontakter som vi har haft under denna tid .
Tillåt mig även att än en gång tacka min medföredragande , Leinen , för allt vårt samarbete .
Herr talman , kära kolleger !
Den regeringskonferens som skall starta är viktig , både rent allmänt , men särskilt med tanke på den förestående utvidgningen .
Vid denna skall den struktur och den metod som skall ligga till grund för Europas funktion i det 21 : a århundradet utarbetas .
För att Europeiska unionen i framtiden skall kunna fungera effektivare , mer demokratiskt och med full öppenhet , är det uppenbart att det krävs en omfattande och grundlig reform av Europeiska unionens institutioner liksom av deras arbetsmetoder .
Av avgörande betydelse för att denna reform skall lyckas är den dagordning som skall ligga till grund för arbetet på regeringskonferensen .
Av besluten från toppmötet i Helsingfors framgår att den dagordning som man där kom överens om inte är tillfredsställande , och att den inte garanterar de nödvändiga och påtagliga förändringar som är ett måste för att skapa ett Europa som fungerar bättre , är effektivare , mer demokratiskt och mer öppet .
Och detta på grund av att den är begränsad till endast de tre frågor som på ett lösryckt sätt berör strukturen och funktionen hos endast två av Europeiska unionens institutioner .
Jag skall inte upprepa det , för ni känner väl till det allihop .
Detta mitt konstaterande berättigas dels av det ständiga kravet från de europeiska medborgarna , som till och från är mycket kraftigt , dels av de enorma dimensionerna på det projekt som Europeiska unionen redan har gett sig in i , utvidgningen .
Mot denna bakgrund är det inte möjligt att man i dagordningen för den nya regeringskonferensen inte inbegriper frågor som , om de får en lösning , skulle säkerställa en smidig funktion för alla - inte bara vissa - av Europeiska unionens institutioner .
Liksom det inte heller är möjligt att man i dagordningen inte inbegriper frågor som dagligen berör och som därför är mycket påtagliga för den europeiska medborgaren .
Herr talman , kära kolleger !
Europaparlamentet har under sina många diskussioner och i de betänkanden som har lagts fram till dags dato öppet varit för att sammankalla en regeringskonferens .
Jag begär emellertid att man på denna parallellt skall ta upp både frågor som förbättrar och fullbordar reformen av - och jag upprepar det - alla institutioner och frågor som direkt berör och intresserar de europeiska medborgarna .
Som till exempel hälsa , energi , kultur , transport och till och med turism .
Vad gäller frågan om dagordningen till slut kommer att utvidgas eller inte , är den å ena sidan fortfarande under diskussion .
Och här vill jag verkligen prisa det sätt på vilket det portugisiska ordförandeskapet , som vid upprepade tillfällen inför Europaparlamentet har förbundit sig att arbeta i den riktningen , har uppträtt politiskt .
Å andra sidan får en ökning eller ett bevarande av antalet frågor inte under några omständigheter leda till att den betydelse som varje medlemsland tillskriver regeringskonferensen minskar .
Och detta av den anledningen att den institutionella ram som skall ligga till grund för Europa i framtiden är en grundläggande princip för den europeiska integreringen och följaktligen en fråga av högsta nationella betydelse för varje land som är medlem i unionen .
Herr talman , kära kolleger !
Med detta som bakgrund uppmanar jag kammaren att godkänna det yttrande som jag och Leinen har lagt fram , så att regeringskonferensens arbete kan komma igång den 14 februari och så att våra två företrädare på denna , Brok och Tsatsos , kan gå framåt med Europaparlamentets samtycke i det svåra arbete som de har framför sig .
Samma sak gäller även för Europeiska kommissionen , och jag vill , återigen , tacka kommissionär Barnier för hans kontakter med Europaparlamentet och för de mycket konstruktiva förslag som han har lagt fram för oss .
Herr talman , herr rådsordförande , herr kommissionär !
Jag är ense med min medföredragande Dimitrakopoulos om att den dagordning man beslutade om i Helsingfors inte räcker till för att behärska de utmaningar som en utvidgning med 13 nya stater innebär .
Enligt vår åsikt skulle en minireform innebära att vi går miste om en chans .
Minireformen skulle också äventyra Europeiska unionens stabilitet .
Att Europeiska unionen på så vis skulle äventyras genom att den tänjs ut för mycket och fördjupas för litet kan och får Europaparlamentet inte acceptera .
Vi vill här än en gång erinra regeringarna om att parlamentet måste ge sitt godkännande innan en ny medlem tas upp i unionen .
Detta beslut om utvidgningen kommer parlamentet säkerligen också att fatta i ljuset av resultaten från denna regeringskonferens .
Vi fastslog den 18 november 1999 hörnstenarna i vår dagordning för denna regeringskonferens 2000 .
Jag vill bara än en gång nämna några punkter : Föreskrifter för ett förstärkt samarbete med dessa 20 och 25 medlemsländer , integrationen av säkerhets- och försvarspolitiken inom gemenskapens ram , införlivandet av stadgan för de medborgerliga rättigheterna i det nya fördraget , en konstitutionalisering av unionen genom att man delar upp fördragen i en grundläggande del och en andra del , reformen av artikel 48 , så att parlamentet vid kommande ändringar i fördraget också faktiskt får delta jämställt vid sådana förhandlingar , och - det vill jag också nämna - en stadga för europeiska partier , så att nästa Europaval verkligen gäller europeiska frågor och inte blir någon nationell inrikespolitisk uppgörelse .
Slutligen också stärkandet av institutioner och instrument för gemenskapens ekonomiska och sociala politik samt sysselsättningspolitik som jämvikt till den europeiska integrationen av valutan och de gemensamma pengar , som vi ju redan har beslutat om .
Vid sidan av en utvidgad dagordning vill vi också ha en förbättrad metod för utarbetandet av detta nya Europafördrag .
För medborgarnas skull måste det garanteras en större öppenhet i den politiska processen under regeringskonferensen .
Därför kräver vi ett omfattande deltagande från parlamentets sida på alla nivåer .
Unionen har en dubbel legitimitet , den är en union av stater , men också en union av folk .
Det vore på tiden att detta också finner sitt uttryck i metoden för att utarbeta ett nytt fördrag .
Företrädarna för Europaparlamentet bör då också verkligen delta i den grupp som förbereder det , både på ministernivå och på Europeiska rådets sammanträde , såvitt detta råd ägnar sig åt regeringskonferensen .
Regeringarna har beslutat att öppna denna regeringskonferens den 14 februari .
Parlamentet kommer i morgon under detta minisammanträde att avge sitt yttrande och därigenom skapa förutsättningar för regeringskonferensen att börja .
Jag vill inte dölja att många kolleger hellre skulle ha väntat tills vi fått en rapport från det portugisiska ordförandeskapet efter dess besök i huvudstäderna , för att få veta om det finns någon rörelse eller dynamik för en utvidgad dagordning .
Men vi har förtroende för att det portugisiska ordförandeskapet , med det engagemang som det har visat här , vid toppmötet i mars i Lissabon kommer att föreslå ytterligare punkter för dagordningen .
Vi ber regeringarna att följa detta förslag från det portugisiska ordförandeskapet .
Såtillvida finns det här ett förtroendeförskott , och vi hoppas verkligen att vi inte blir besvikna om vi redan nu avger vårt yttrande utan att exakt känna till vad som nu finns i fråga om ny dynamik och vilka de ytterligare punkterna på agendan kommer att bli .
Det yttrande som vi lägger fram för er är en tydlig signal till regeringarna att inte missa den sista chansen att före utvidgningen genomföra en ambitiös reform av EU och höja acceptansen för detta nästa Europafördrag , där det finns en större öppenhet och där parlamentets fullständiga deltagande garanteras .
Även jag vill tacka det portugisiska ordförandeskapet , och tacka kommissionär Barnier för samarbetet .
Jag ber om stor samstämmighet här i parlamentet för att godkänna vårt yttrande .
Herr talman , ärade kollegor !
Först och främst vill jag tacka föregående två talare för visat förtroende för det portugisiska ordförandeskapets arbete i frågan .
Jag tror att jag från sammanträdet i utskottet för konstitutionella frågor - senare bekräftat av portugisiska utrikesministerns uttalanden under plenarsammanträdet i parlamentet - väl har klargjort att Portugal ser sig själv som den drivande kraften bakom regeringskonferensen .
Vi tror faktiskt att det här är ett ypperligt tillfälle för en utvidgning av unionen , men vi måste handla snabbt så att vår strävan kan kombineras med vårt behov av att nå resultat fram till årets slut .
Det är ett problem som vi alla ställs inför , utan tvivel förstärkt av de svårigheter som en del regeringar har med att få igenom vissa åtgärder i sina parlament eller via eventuella nationella folkomröstningar .
Vi måste komma ihåg att vi står inför en nästan två år lång ratificeringsprocess och att det är viktigt att vi ser till att den blir framgångsrik .
Vilken hypotes som helst om ett misslyckande är ett globalt misslyckande för unionen .
Vi måste därför se till att slutresultatet av konferensarbetet är något så när rimligt och tillräckligt accepterat av allmänheten och ländernas politiska grupperingar .
Våra förslag inför konferensen mottogs enligt min mening mycket väl av de olika regeringarna .
Inrättandet av den förberedande grupp jag själv är ordförande i var också ett svar på Europaparlamentets oro över ledamöternas grad av inblandning i det här läget av förhandlingarna .
Jag räknar därför med våra vänner Brok och Tsatsos arbete , ett arbete som tveklöst kommer att vara till stor nytta i den debatt som skall föras inom gruppen .
Jag vill tillägga att det är vår tolkning som med er medverkan kommer att göras i plenum , precis som vilken annan av en medlemsstat utsedd gruppmedlem eller kommissionsledamot .
Jag menar också att portugisiska ordförandeskapets beslut att utse utrikesministern till ordförande och leda ministergruppen också skall tolkas som att man ville försäkra Europaparlamentets talman om en så jämbördig företrädare som möjligt och inte någon som skulle kunna anses som mindre värdig talmannen i en institution som denna .
Fru talman , ärade kollegor , det är svårt att göra en sammanfattning av de kontakter - och meningen med de kontakter - jag har haft med de olika länderna , jag har ju ännu inte hunnit avsluta min rundtur bland huvudstäderna under vilken jag försökte ta reda på hur länderna ser på konferensen och vilka förväntningarna är .
Jag tror dock att jag avslutningsvis kan säga att flertalet länder verkar vara beredda att inleda debatten , vilket inte nödvändigtvis betyder att man är beredd att avsluta på ett sätt som står i samklang med parlamentets tolkning av vissa nödvändiga reformer , något som vi från och med nu måste ha i åtanke .
Det finns i alla fall en öppning , från flera regeringars sida , såtillvida att man kan acceptera många av de ämnen jag föreslog .
Det är självklart att ämnen av det här slaget hör ihop med frågor av institutionell natur , något som det portugisiska ordförandeskapet menar skall ingå i dess mandat .
Detta vill jag gärna klargöra : Vårt mandat , mandatet som härrör från Helsingfors är inte bara från portugisiskt håll sett ett mandat från de tre left overs från Amsterdam .
Det mandat vi fick med oss från Helsingfors är de tre left overs från Amsterdam , men det rör sig också om institutionella frågor .
Här har vi givetvis det arbete som kan associeras med gemenskapsinstitutionerna , unionens myndigheter , problemet med ett förstärkt samarbete , en fråga som kan förknippas med alla left overs i ordets egentliga bemärkelse , men även med frågor som exempelvis unionens juridiska karaktär , förenklingen av fördragen liksom andra frågor som på ett organiskt sätt har att göra med en revision av Fördraget om Europeiska unionen och som vi menar är viktiga , nämligen de som har att göra med parlamentets struktur vid en utvidgning i efterhand , de övergångsbestämmelser som måste verkställas om utvidgning sker före utgången av parlamentets mandatperiod , liksom kommissionärernas personliga ansvar .
Nåväl , en rad frågor som vi menar att vi kan och bör sätta upp på konferensens dagordning .
Från medlemsstaternas sida har vi sett en antydan till att kunna acceptera en sådan möjlighet .
Jag vill säga att min avsikt är att initiativen under det portugisiska ordförandeskapet snabbt och med påtaglig grund skall inledas och sättas igång .
Jag har inte för avsikt att lansera de förberedande gruppernas arbeten som en enkel liten ämnesgranskning , en slags notarie som står på flera medlemsländers sida .
Jag tänker inte utge mig för att vara en notarie , jag tänker lägga fram konkreta förslag angående vissa frågor , där jag givetvis löper risken att förslagen inte får ett gott mottagande .
Vår avsikt är att dela upp den förberedande gruppens arbete i två perioder under vilka alla ämnen kommer att analyseras .
Den första perioden kommer att inledas med en omröstning med kvalificerad majoritet , därefter försöker vi identifiera de institutionella frågor som har att göra med left overs , och först därefter tar vi itu med frågan om kommissionen och röstfunderingarna .
Det förstärkta samarbetet kommer att tas upp i samband med de institutionella frågorna .
Avslutningsvis , under andra perioden , tänkte vi än en gång titta på de frågor som under tiden redan har behandlats , som har granskats vid ministersammanträdena , samt titta på de frågor som uppstått allt efter arbetets gång .
Här är det viktigt att veta om institutionernas diskussionen om säkerhets- och försvarsfrågor har mognat så att vi kan inkludera dem i slutfasen av konferensen .
Detsamma kan sägas om dokumentet om de grundläggande rättigheterna .
Vi får se om den debatt som skall föras vid institutionerna om den här frågan kan få oss att dra den slutsatsen att ta med den i regeringskonferensen , det vill säga under årets andra hälft .
Detta är i princip ordförandeskapets avsikt .
Vi kommer att avge en rapport till Europeiska rådet i Lissabon , en rapport som givetvis måste baseras på sakuppgifter , eftersom rapporten skrivs i mars och konferensen bara började i februari .
Vi hoppas att den andra rapporten , den rapport som ordförandeskapet kommer att lämna vid det andra Europeiska rådet , kommer att vara mera substantiell och något mera konkret , konkret när det gäller fördragstexterna , om nu det är möjligt .
Vi noterar kommissionens förslag .
Ordförandeskapet kommer att ta emot förslagen och på lämpligt sätt ta upp dem till behandling under konferensen , oberoende av detta kan varje medlemsstat begrunda de lösningar som kommissionen föregriper i sitt förslag .
Vi hoppas kunna inkludera alla förslag och dokument som medlemsstaterna kan tänkas skicka oss i den här frågan .
För övrigt kommer vi att vädja till medlemsländerna att så fort som möjligt sända in sina bidrag till konferensen så att de inte ankommer för sent .
Konferensen är alltid öppen för förslag från medlemsländerna , men vi vill att de snarast definierar sina ståndpunkter .
Fru talman och ärade kollegor , detta är enligt vår mening det viktiga med konferensen .
Från vår sida är vi med andra ord fast beslutna att arbetet under halvåret med portugisiskt ordförandeskap , under vilket regeringskonferensen äger rum , blir effektivt och seriöst .
Vi hoppas att vi till det franska ordförandeskapet kan överlämna något påtagligt och i viss mån representativt för de tendenser som har sprungit fram hos medlemsländerna under arbetets gång .
Herr talman !
Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater var inte nöjda med resultatet från Europeiska rådets möte i Helsingfors .
Vi ansåg att dagordningen var för begränsad , för vår grupp utgick från fördragets logik , närmare bestämt från protokollet om unionens institutioner .
I Helsingfors kom regeringarna överens om att en minimireform är tillräcklig , så länge Europeiska unionen består av mindre än 21 stater ; dessutom krävs det en djupgående reform .
Samtidigt godkände Europeiska rådet i Helsingfors en utvidgning med 13 nya medlemsstater .
Det finns således en motsägelse i att påbörja anslutningsförhandlingarna med 13 samtidigt som man vill ha en minimireform .
Vi tillämpar fördragets logik och vill att dagordningen för nästa regeringskonferens skall rymma en mer djupgående reform av unionen .
Det är anledningen , herr talman , till att vi håller denna debatt i parlamentet i dag , eftersom vi inte vill skjuta upp inledandet av konferensen .
Rent teoretiskt hade vi kunnat göra det .
Vi hade kunnat rösta den sjuttonde den här månaden , och då hade inte konferensen kunnat börja den fjortonde .
Men det ville vi inte göra , för vi vill ge regeringarna och kandidatländerna en tydlig politisk signal om att vi önskar genomdriva denna reform just för att underlätta en utvidgning .
Herr talman , jag är glad över att kunna framföra detta till det portugisiska ordförandeskapet , för de har vunnit ett gott anseende här i parlamentet .
Det portugisiska ordförandeskapet delar många av parlamentets ambitioner , och man har lovat att göra vad man kan för att regeringskonferensens dagordning skall fyllas på med andra frågor som är av största vikt .
Och jag vill dessutom påpeka , herr talman , att Europaparlamentets ambitioner inte är ambitioner för parlamentets egen räkning .
Europaparlamentet kommer hur som helst att stärkas politiskt av det fördrag som regeringskonferensen resulterar i .
Anledningen till detta är mycket enkel : Under regeringskonferensen kommer man , i enlighet med överenskommelsen i Helsingfors , att ta ställning till vilka av de frågor som hittills har avgjorts med enhällighet som skall avgöras med kvalificerad majoritet .
Det innebär att antalet frågor som avgörs med kvalificerad majoritet kommer att öka .
Och det framgår redan av gemenskapens regelverk att de lagstiftningsfrågor som avgörs med kvalificerad majoritet även skall vara föremål för parlamentets medbeslutande .
Därför innebär en ökning av den kvalificerade majoriteten en ökning av parlamentets medbeslutande .
Däremot skulle parlamentet inte uppfylla sin roll som en supranationell europeisk institution om det inte tänkte på unionens politiska utformning .
Det är det vi ägnar oss åt nu .
Vi anser att unionens politiska utformning förutsätter att även andra frågor behandlas .
Bland annat sådana som handlar om införandet i fördraget av säkerhets- och försvarsfrågor , frågor vars betydelse har ökat markant den senaste tiden och därför bör införlivas i fördraget .
Förvisso även stadgan om de grundläggande rättigheterna i Europeiska unionen , vars utformning påbörjades i går , och jag tror att man gripit sig an den uppgiften på ett mycket positivt sätt .
Vi kommer i stor utsträckning att verka för att européerna skall bli medvetna om fördelarna med att vara europé och att en europeisk medborgare har vissa grundläggande rättigheter som är knutna till unionens institutioner .
De förslag , herr talman , som vi konkretiserar i ett annat betänkande , utgör tillsammans med kommissionens förslag ett utmärkt dokument som - vilket jag nu har nöjet att få säga till herr Barnier - således kommer att vara ett underlag till regeringskonferensen .
Det får vi tala mer om en annan dag .
I dag måste vi ge klartecken till sammankallandet av denna konferens , och Europeiska folkpartiets grupp , herr talman , är beredd att ge klartecken .
Herr talman !
Å socialistgruppens vägnar kan jag framföra att vi kommer att stödja det förslag till yttrande som lagts fram av föredragandena för utskottet för konstitutionella frågor .
Vi avger ett positivt yttrande om att sammankalla regeringskonferensen helt enkelt därför att vi är mycket imponerade av det portugisiska ordförandeskapet som har gått med på vår begäran om att dagordningen för regeringskonferensen utvidgas .
Resterna från Amsterdam är inte ett bra uttryck eftersom de är mycket viktiga frågor i sig själva .
Låt oss kalla dem de tre första punkterna för regeringskonferensen .
Dessa tre första punkter är mycket viktiga , men detta är frågor som diskuterades noga av våra medlemsstater under den senaste regeringskonferensen .
De kom inte helt fram till en slutsats om dem men det krävs verkligen inte nio månader av ytterligare granskning av dem .
De kräver en politisk överenskommelse .
Det är mer en fråga om nio minuter , kanske nio timmar om det är svårlöst , inlåsta tillsammans i ett rum för att nå en lösning om dessa frågor , inte nio månader .
Under dessa omständigheter skulle det vara dumt att inte utvidga dagordningen .
Det finns andra frågor som borde vara givande att granska framför allt före en så stor utvidgning av unionen med så många nya länder .
Ingen begär att det ska vara julklappsstämning .
Ingen begär en regeringskonferens i stil med Maastricht med hundra eller fler punkter att diskutera .
Men det finns sex , sju , åtta , kanske nio punkter som det skulle vara mycket lämpligt och nyttigt att få en lösning på .
Det finns tid .
Kom ihåg regeringskonferensen som ledde fram till Europeiska enhetsakten .
Den pågick bara fem månader .
Den regeringskonferens som ledde fram till det enorma Maastrichtfördraget pågick ett år .
Enbart konferensen om Amsterdamfördraget pågick i ett och ett halvt år och det berodde på att alla visste att man måste vänta på resultaten av det brittiska valet om man skulle få något resultat från den regeringskonferensen , så det var av en annan orsak .
Ett år är tillräcklig tid för att lösa en stort antal frågor , och det borde utan tvivel vara tillräcklig tid för att lösa de få avgörande frågor som vi önskar lägga till på dagordningen .
Jag är glad att kommissionen delar vår åsikt .
Kommissionen har just offentliggjort sitt yttrande och den har gjort exakt det som parlamentet begärde av den - att lägga fram ett fullständigt och samlat förslag med verkliga förslag till fördragsartiklar .
Jag tackar kommissionen för detta även om jag naturligtvis inte är överens med allt det som kommissionen framförde .
Jag anser att det finns några brister i det som den presenterade .
Hur som helst har kommissionen tillhandahållit en tjänst och jag uppskattar att kommissionär Barnier som finns här bland oss i dag för att han gjorde detta .
Den har för allmänheten presenterat några av de avgörande frågor som vi måste lösa under denna regeringskonferens .
Det är alltsammans bara bra .
Parlamentet , rådets ordförandeskap och kommissionen drar åt samma håll för att få en bredare dagordning .
Jag önskar er all framgång , rådets ordförande , för att se till att Europeiska rådet godkänner denna dagordning och att på Alla hjärtans dag när ni inleder regeringskonferensen det kommer att ske under gynnsamma omständigheter och att ni kommer att kunna slutföra den på ett bra sätt , även när det franska ordförandeskapet tar över i slutet av detta år .
Vi skall inte längre oroa oss över att dagordningen för regeringskonferensen skall bli begränsad .
Det är en av de politiska slutsatserna som vi måste dra från det allvarliga beslutet av 14 medlemsstater i går att i verkligheten frysa våra förbindelser med en partner .
Det gör det omöjligt för dessa samma medlemsstater att vid regeringskonferensen misslyckas med att ge en effektiv mening vad gäller skydd och främjande av grundläggande fri- och rättigheter .
Det är redan konstigt att inom det konvent som tar fram förslag till stadgan se företrädare från några medlemsstater , särskilt Storbritannien och Frankrike , försöka argumentera att en obligatorisk stadga på något sätt skulle vara en kränkning av nationellt självbestämmande .
Det är viktigt att regeringskonferensen förbereder hur införandet av en ordning för grundläggande fri- och rättigheter inom fördraget godkänns .
En del av detta är att förbättra medborgarnas möjlighet att väcka talan vid domstol .
Ett annat sätt är att själva unionen undertecknar Europakonventionen .
Ett annat sätt är utan tvivel att nationella parlament och nationella politiska partier finna en kraftfullare roll som de kan spela inom Europeiska unionens verksamhet och att dela ansvaret för att skapa europeisk parlamentarisk demokrati .
Min grupp välkomnar absolut regeringskonferensen och kommer att medverka i denna fördragsreform i största möjliga grad .
Herr talman !
Gruppen De Gröna / Europeiska fria alliansen anser att Europaparlamentets beslut att skyndsamt yttra sig om regeringskonferensen neutraliserar den politiska betydelsen av uppmaningen till rådet och gör den , i slutändan , ganska ointressant .
Vi hade hellre velat få en tydligare uppfattning om dagordningen , något större säkerhet vad gäller metoden , innan vi avger vårt yttrande , och vi uppskattar inte den bristande respekt som det portugisiska ordförandeskapet visade Europaparlamentet genom att bestämma att regeringskonferensen skulle börja på Alla hjärtans dag , den första dagen under sammanträdesperioden i Strasbourg .
Jag tror dessutom att eftersom detta är ett ganska viktigt yttrande , så kan vi också rösta för det och jag tror att majoriteten i vår grupp kommer att rösta för det .
Man jag vill ändå understryka att det är ganska grymt att se hur litet intresse denna reform väcker .
Händelserna i Österrike visar på ett mycket tydligt sätt behovet av en reform , en struktur för den europeiska demokratin , för att bestämma de principer som samtliga medlemsstater skall ansluta sig till .
Det smärtar också att tänka sig att initiativet gentemot Österrike i verkligheten är frukten av en överenskommelse mellan regeringar och att Europeiska unionen och dess institutioner inte hade möjligheter eller den gemensamma kraften att agera för att förhindra utvecklingen och leda in den på andra banor .
Jag tror att detta är något som vi måste reagera mot , detta måste vi göra under regeringskonferensen och jag hoppas verkligen att Europaparlamentet inte med det här yttrandet , som avgivits med sådan ovilja , helt har uttömt sin förmåga att utöva påtryckningar på rådet och medlemsstaterna för att denna regeringskonferens inte bara skall bli en rent teknisk övning utan väcker den entusiasm som vi fick se spår av i detta parlament för några timmar sedan .
Herr talman , herr rådsordförande , herr kommissionär , ärade kolleger !
Jag anser att man inte tillräckligt ofta och ljudligt kan säga att den föredragningslista som rådet har fastställt för regeringskonferensen är politiskt fullständigt oacceptabel , och jag vill tillfoga att jag anser att den rent av är skamlig .
Vi befinner oss nämligen i en historisk situation , där man förhandlar respektive kommer att ta upp förhandlingar med 12 stater , och nu befinner vi oss gemensamt i en situation där det inom överskådlig tid kan bli verklighet att Europa växer samman .
Men hur skall då unionen kunna utvidgas , om man inte nu - alltså före utvidgningen - ser till att man har effektiva verktyg ?
Därför är vi som grupp positiva till regeringskonferensen .
Vi anser att den är absolut nödvändig och brådskande och vi hoppas att den i själva verket skall åstadkomma resultat som möjliggör en snar utvidgning av Europeiska unionen .
Min grupp , herr rådsordförande , har med tillfredsställelse noterat att rådets ordförandeskap inte är tillfreds med den nuvarande situationen .
Därför kan ni vara säkra på att även Gruppen Europeiska enade vänstern / Nordisk grön vänster kommer att arbeta för att unionen äntligen skall göra sina hemläxor .
Det handlar om varken mer eller mindre än Europas framtid , och det handlar framför allt om ett Europa som medborgarna faktiskt uppfattar som sitt eget , eftersom de kan vara med och utforma det , och eftersom de bekymmer och trångmål , problem och frågor som de dagligen möter också tas på allvar i politiken .
De slutna dörrarnas politik , samråden i den stilla kammaren , allt detta måste en gång för alla förpassas till det förflutna .
Därför krävs det öppenhet .
Jag anser att ni som ordförandeskap bör se till att tåget inte fortsätter att gå som hittills , och att människorna inte blir stående kvar på perrongen som fördragsanalfabeter .
Vi anser att det är absolut nödvändigt att man inte bara gör allt för att ge medborgarna omfattande information om vad som sker vid regeringskonferensen och resultaten av den , utan de måste snarare integreras direkt i hela reformprocessen .
Vi anser också att de politiska beslutsfattarna äntligen måste hoppa över sin skugga och efter regeringskonferensen fråga medborgarna i folkomröstningar om de är införstådda med hur deras Europa kommer att utvecklas i framtiden .
På så vis skulle vi faktiskt få ett medborgarnas Europa , och vi skulle faktiskt få en helt ny kvalitet med demokratisk legitimitet för unionen .
Jag vill klart och tydligt ta upp en annan central demokratifråga .
Som ledamot av den församling , som nu har påbörjat sitt arbete på stadgan för de grundläggande rättigheterna , vill jag klart säga : För mig och min grupp räcker det inte med att högtidligt förkunna stadgan .
Vad kommer väl medborgarna att säga när man högtidligt förkunnar rättigheter för dem , medan de inte som individer kan överklaga något ?
Nej , jag tror att det bara skulle fördjupa unionens trovärdighetskris ännu mer .
Det dåliga valdeltagandet vid Europavalen bör verkligen vara en tillräcklig larmsignal för alla .
Det vi behöver är synliga rättigheter för var och en , stadgan om de grundläggande rättigheterna måste blir bindande rätt för alla människor som bor i unionen , för alla dess medborgare .
Detta är det mål som vi för medborgarnas skull gemensamt bör arbeta för , och jag förväntar mig av regeringskonferensen att beslutet från Köln i denna fråga revideras vid årets slut .
Naturligtvis handlar det också om att man har effektiva beslut och fungerande institutioner i en union med 27 och fler medlemsstater .
Med enbart en liten minireform , som rådet har bestämt sig för , kommer det inte att lyckas , och därför bör alla institutioner prövas .
Vi behöver modiga förändringar , och därvid måste vi samtidigt se till att man ägnar största uppmärksamhet åt jämställdheten mellan de stora och de små staterna .
Detta vill jag särskilt betona som ledamot från ett stort medlemsland .
Jag tackar kommissionen för de förslag den har lagt fram , och jag är säker på att vi här kommer att få omfattande diskussioner med medborgarna även i Europaparlamentet om alla de frågor som de har framkastat .
Jag vill också ta upp en sista fråga .
I parlamentets yttrande krävs det uttryckligen ändringar av fördraget när det gäller den ekonomiska politiken .
I själva verket är det så att globaliseringen av samhällsekonomin , men framför allt införandet av euron och den stabilitetspakt som är förbunden därmed , gör det nödvändigt att inte bara fråga efter bakgrunden till beslutsprocesserna .
Det som framför allt krävs är modet att kritiskt granska unionens hittillsvarande politik .
Det handlar om ett socialt rättvist Europa .
Ett socialt rättvist Europa är oförändrat högaktuellt , ty det handlar i första hand om att målinriktat ställa kampen mot massarbetslösheten och fattigdomen i centrum för unionens politik .
Hit hör därför också , enligt min åsikt , modet att ändra artikel 4 i EG-fördraget , som unionen på klassiskt nyliberalt vis definierar som en öppen marknadsekonomi med fri konkurrens , och dit hör enligt min åsikt även artikel 105 i EG-fördraget , ty Europeiska centralbanken måste äntligen få ett i fördraget fastslaget politiskt uppdrag att med sin penningpolitik främja hållbar tillväxt och sysselsättning .
Herr talman !
Gruppen Unionen för nationernas Europa anser att dagordningen för nästa regeringskonferens , såsom den fastställts av Europeiska rådet i Helsingfors , dvs. strikt inriktad på frågor om beslutsfattande i ett utvidgat Europa , måste respekteras .
Den måste respekteras med tanke på att konferensen behöver utföra ett effektivt och snabbt arbete före utvidgningen .
Det är anledningen till att vi inte kan ansluta oss vare sig till Europaparlamentets ståndpunkt eller till kommissionens , som alltför mycket vill utvidga denna dagordning och dessutom utvidga den i fel riktning , dvs. i riktning mot en centralisering och en allt hårdare låsning av det europeiska systemet.Vår grupp har därför lämnat in en rad ändringsförslag som , i tur och ordning , bildar en verklig alternativ resolution .
Vi säger där att nästa regeringskonferens måste överväga ett beslutssystem som bättre respekterar den nationella suveräniteten .
Vi beklagar att kommissionen i sitt yttrande av den 26 januari envisas med att fortsätta rutinvägen med ett likriktat Europa utvidgat mot öster , en centraliserad superstat som fungerar med hjälp av majoritetsbeslut .
Federalisterna tror att de på så sätt skall kunna skapa enhet genom tvång , men det är en fullständigt ytlig idé .
Tvärtom , herr talman !
I ett utvidgat Europa kan likriktningen som påtvingas genom ett felaktigt användande av majoritetsbeslut bara leda till explosion .
Det europeiska centraliserade systemet , såsom det utvecklas i dag och så som vi kan extrapolera det , pressar samman nationerna och därigenom pressas också den nationella patriotismen samman , den som utgör hjärtat i vår försvarsvilja .
Det Europa som då uppstår är inte starkare utan svagare , eftersom det inte vet vem det är eller vad det försvarar .
Det är anledningen till att vi alltid sagt att utvidgningen bara är möjlig genom att vi klart accepterar mångfalden och friheten för de folk som utgör Europa , dvs. genom att anta en variabel geometri som bygger på respekt för den nationella självständigheten .
Vi gläds i dag åt att se att denna idé gör framsteg i miljöer som tyvärr fortfarande ligger utanför Europaparlamentet och kommissionen.Ett Europa med variabel geometri är ett Europa som respekterar sina nationella demokratier , som stöder sig på sina nationer , på sin nationella patriotism , i stället för att hela tiden förfölja dem .
Det är där vi hämtar viljan att försvara oss mot yttre hot och inte beslutsförfaranden som är tvingande och konstlade och som kommissionen fått för sig att föreslå den kommande regeringskonferensen .
Herr talman , kära kolleger !
Jag talar som företrädare för de italienska radikala ledamöterna och jag skulle vilja säga till rådets ordförande att han förmodligen har kunnat konstatera vad som är parlamentets uppgift .
Det är knappast en slump att det sista inlägget var det enda som han instämde i helhjärtat - jag säger detta utan att på minsta sätt ironisera över den position , som är fullständigt respektabel , som Berthu och hans grupp har intagit - men det är ingen slump att Europeiska rådets beslut stöds av dem som egentligen befinner sig i detta parlament enbart för att de är motståndare till - något som är fullständigt respektabelt - en ytterligare integration i Europa .
Detta är det budskap som parlamentet skickar till rådet .
Jag hoppas att det portugisiska ordförandeskapet - och som även jag vill gratulera - kan överbringa detta parlaments budskap och blir de som bär fram resultatet av vårt kompromissarbete till St. Valentins altare , men under alla omständigheter kommer vi i morgon att yttra oss negativt om dagordningen för regeringskonferensen .
Det här budskapet måste bli mycket tydligt : det är så vi tolkar den röst som vi avger i morgon .
Vi avger ett yttrande - som är tekniskt och juridiskt nödvändigt - för att sammankalla regeringskonferensen den 14 februari , men vi yttrar oss negativt om innehållet .
Det räcker att betänka de faktiska omständigheterna : vi såg Österrike för ett tag sedan , men vi kan också se på aktiebörserna , herr talman : när , på ett år , det stora europrojektet kan förlora 16 procent gentemot dollarn så borde kanske inte en regering , men väl en god familjefader , fråga sig om man kan säga till medborgarna att det enda man kan förhandla om är antalet europeiska kommissionärer eller andra frågor av samma typ .
Det är uppenbart att målet måste vara ambitiösare .
Vi radikala har lagt fram ändringsförslag som vi kommer att underställa kammaren , för att skärpa texten , för att till exempel begära det som borde vara ett minimum - om man nu skall tala om artikel 6 och 7 - dvs. att den europeiska konstitutionen även skall utformas av Europaparlamentet , att man föreslår att ändringarna i fördraget skall godkännas av Europaparlamentet .
Vi vet att det även finns andra frågor : till exempel har många kolleger , tillsammans med oss , skrivit under frågan om var institutionerna skall vara belägna , en fråga som vi tycker borde utgöra en del av de diskussioner som förs under regeringskonferensen .
Låt mig avslutningsvis hoppas att det budskap som vi ger i morgon blir ett kraftfullt budskap , för en gångs skull betydelsefullt , och att man verkligen , även tack vare de ansträngningar som det portugisiska ordförandeskapet gjort , kan revidera denna dagordning , för annars tror jag verkligen att detta är ett tillfälle som går förlorat , inte bara för ögonblicket , utan för många år framåt .
Herr talman !
Kommissionens ordförande var inte helt ärlig när han i förra veckan uttalade sig om regeringskonferensen .
Han sade att det fortfarande skulle finnas enhällighet i sociala frågor , men i kommissionens förslag vill man ju uttryckligen ha majoritetsbeslut i socialförsäkringsfrågor och frågor som rör de skatter som har samband med den inre marknaden , och det betyder att huvuddelen av de sociala systemen i medlemsstaterna skall kunna ändras av en majoritet i Bryssel , även om en enhällig fransk nationalförsamling , ett enhälligt brittiskt underhus och en enhällig nederländsk andrakammare är emot det .
Man går här in i folkstyrets hjärta rörande fördelningspolitiken och medborgarnas sociala villkor , som är det man vill påverka när man går till val .
Detta skall vi inte längre kunna bestämma över som väljare .
Detta skall vi inte längre kunna ändra på valdagen .
Bryssel vet bättre .
Prodi bebådade också större öppenhet , men hans förslag till förordning innebär en direkt bakåtsträvande utveckling och det är inte bara min , utan också Europeiska ombudsmannens uppfattning .
I dag är kommissionen skyldig att individuellt väga sekretesshänsynen mot medborgarnas krav och förväntningar rörande öppenhet , och om kommissionens förordning antas kommer kommissionen att ha att utestänga en rad dokumentkategorier , utan att genomföra en konkret bedömning .
Man vill också skapa rättsliga krav på sekretess och sekretessbelägga dokument som i dag är offentliga i en rad medlemsstater .
Under titeln " utveckling för öppenhet " gör man att en rad dokument inte blir tillgängliga för allmänheten .
Det är mycket orwellskt .
Jag vill be Prodi att aldrig mer kommentera ett förslag här i kammaren , som inte samtidigt finns tillgängligt för allmänhetens kritiska kontroll .
Prodi talade i positiva ordalag om ett förslag som annars hade fått kritik , då det i det nya förslaget till förordning framställs som ett framsteg att man nu skall skapa insyn i alla dokument som finns hos kommissionen , men efteråt kommer en lång , lång lista över undantag , och det finns rättsliga krav på sekretess rörande dessa undantag .
I den franska texten står det " refuse " , i den engelska " shall " , vilket innebär att kommissionen skall hemlighålla uppgifter som i dag är offentliga i t.ex. mitt hemland .
Det finns också en gummiparagraf om förhandlingarnas och institutionernas effektivitet , som kan användas till vad som helst , det är därför ...
( Talmannen avbryter talaren . ) .
Herr talman , kolleger !
Efter det portugisiska ordförandeskapets framställning har jag en känsla av att man tar itu med denna regeringskonferens med väl övervägda tankar och ett stort mått av öppenhet .
Som Europaparlament kommer vi att utnyttja dessa möjligheter för att där på lämpligt sätt lägga fram våra frågor .
Kommissionens hittillsvarande förberedelser går åt rätt håll , även om de också enligt Europaparlamentets resolutioner inte går tillräckligt långt .
Det kommer ju också att diskuteras senare .
Det som är avgörande för denna regeringskonferens är att det uppnås en treklang , nämligen handlingsförmåga , demokratisk legitimitet och öppenhet .
Endast om dessa tre saker finns för handen , får vi till slut en acceptans från medborgarna .
Handlingskraften skall naturligtvis skapas för att det skall vara möjligt för Europeiska unionen att utvidgas .
När vi i denna kammare i dag tidigare förde en annan debatt , så är det ett viktigt tecken för detta .
Vi måste också vara handlingskraftiga i en europeisk union , om det någon gång skulle hända att en regering skulle utöva en totalblockad .
Det är ett viktigt tecken på att majoritetsbeslutet är en avgörande förutsättning för att Europeiska unionen skall kunna arbeta i alla sammanhang .
Detta är särskilt viktigt i samband med utvidgningen , när det gäller lagstiftning , och när det gäller fördrag som för med sig ändringar av lagstiftningen .
Här vill vi naturligtvis också bygga ut motsvarande rättigheter för Europaparlamentet .
Därvid kommer vi som Europaparlament också att agera när det gäller EMU , ty på detta område finns det inte någon tillräcklig kontroll .
Finansministrarna uppträder i Ekofin-rådet och med de 11 staterna i Euro-rådet som om det vore ett evenemang mellan regeringar , vilket inte är acceptabelt .
I motsats till Kaufmann är jag inte positiv till att utvidga kontrollen av Europeiska centralbanken , eftersom jag är för Europeiska centralbankens oberoende .
Men politiskt sett måste kontrollen åstadkommas på lämpligt sätt .
Det gäller också att återställa trojkan kommissionen , rådet och parlamentet i fråga om utrikes- och säkerhetspolitiken , där hittills allt har skötts alltför mycket av rådet , och särskilt de primitiva krisstyrningsåtgärderna , där ansvaret ligger enbart hos kommissionen .
Allt detta har inte tagits med i detta helhetskoncept i tillräcklig omfattning .
Vi måste granska om det är nödvändigt med ändringar här inom ramen för regeringskonferensen .
Rådets portugisiska ordförandeskap har sagt ja till att arrangera överläggningar om detta , för att möjligen få en utvidgning av mandatet .
Jag vill också hänvisa till en annan viktig punkt .
De diskussioner vi i dessa dagar för om exempelvis en regering i ett land i Europa , visar ändå att vi måste fastslå Europeiska unionens intellektuella , moraliska , rättsstatliga inriktning med en gemenskaps- och allmännyttig orientering , och att rättsligt bindande grundläggande rättigheter även av den anledningen måste införas i fördraget , eftersom detta kommer att vara en avgörande stabiliserande faktor .
Jag ber dem som i detta avseende hittills har varit mycket återhållsamma , att överväga om det nu inte är rätt ögonblick att också inse detta sammanhang och kanske ha det mod som krävs , så att vi på lämpligt sätt kan komma vidare med de grundläggande rättigheterna .
Europeiska unionen behöver knappast några nya instrument , inga nya befogenheter .
Det den behöver är instrument för att kunna utnyttja sina befogenheter .
Av den anledningen måste vi se till att instrumenten kan fungera så att vi i medborgarnas namn kan utföra de uppgifter , som vi formellt redan har ålagts i fördraget .
Jag tror att denna regeringskonferens särskilt bör koncentrera sina ansträngningar på detta .
Om vi lyckas uppnå några framsteg här , då kan vi också se fram emot den historiska uppgiften att utvidga Europeiska unionen .
Det måste vara den avgörande punkten .
Ärade ordförandeskap i rådet , jag är övertygad om att det kommer att utformas på ett positivt sätt under er ledning .
Herr rådsordförande !
Ni har säkert , efter att ha lyssnat på de olika inläggen förstått hur uppfattningen att vi skall visa det portugisiska ordförandeskapet förtroende , att vi inte skall öka dess svårigheter genom att skjuta regeringskonferensen på framtiden , har segrat i utskottet för konstitutionella frågor , och även när det gäller ordförandena för de olika politiska grupperna i parlamentet .
Jag kan försäkra er att det inte var lätt att lyckas med detta i förra veckan i det utskott som jag leder , men vi har nu definitivt beslutat att satsa på det portugisiska ordförandeskapet , och det är en satsning som vi verkligen hoppas kommer att gå hem .
Ni talade om era resor mellan olika huvudstäder och ni berättade om de svårigheter som vissa regeringar har att skapa enighet i sina länder och därmed också i sina respektive parlament .
Låt mig påpeka för er att i går genomförde vi en som jag tycker mycket intressant diskussion och dialog med företrädarna för de 15 olika nationella parlamenten , som var närvarande med kvalificerade och engagerade delegationer .
Det handlade inte om att komma fram till några slutsatser - det var inte möjligt att dra några sådana - men diskussionerna var utan tvekan mycket uppmuntrande .
Jag anser att vi måste vara försiktiga , och verkligen vara övertygade om att de olika nationella regeringarna faktiskt försöker övertala sina respektive parlament att ratificera lösningar som motsvarar behovet att utöka unionen och att inte ta skydd bakom motståndet från sina respektive parlament för att inte underteckna de slutsatser som krävs vid regeringskonferensen .
Vi kommer under alla omständigheter att förstärka vårt samarbete , vår dialog med de nationella parlamenten under hela den tid som regeringskonferensen pågår .
I går diskuterade man även inom kommissionen - här företrädd av kommissionär Barnier - som också avgav sitt yttrande .
Man uppskattade ansträngningarna även om man , när det gäller förslagen , uttryckte avvikande åsikter , i likhet med vad även ni har gjort , herr rådsordförande , om jag inte misstar mig .
Det som måste understrykas är det faktum att även i går var många medvetna om risken att utvidgningen leder till att den ursprungliga idén att bygga upp ett politiskt Europa kan komma att ifrågasättas , en risk som för övrigt påpekades i en intervju som inte kan ha undgått någon på grund av den intervjuades auktoritet , nämligen Jacques Delors .
Vi måste därför se till att man vid regeringskonferensen verkligen diskuterar hur man skall förstärka unionens demokratiska bas , hur man skall förstärka - och det har vi redan diskuterat i denna kammare , i samband med situationen i Österrike - systemet av principer , värderingar , rättigheter som ligger till grund för unionen , den roll som de politiska institutionerna skall spela inom unionen , även när det gäller att styra ekonomin .
Vi litar på det portugisiska ordförandeskapet , vi litar på oss själva och vi litar på kommissionen , för allt detta kan man diskutera på ett konstruktivt och produktivt sätt under regeringskonferensen .
Herr talman !
Endast ett förstärkt Europa kommer att klara utvidgningen .
Endast ett förstärkt Europa är osårbart för politiska opportunister som använder sig av ofred .
Därför behövs det grundliga reformer och alltså en utvidgad dagordning för regeringskonferensen .
Det finska ordförandeskapet lyssnade endast till minimalistiska regeringar och var tyvärr stendövt för det här parlamentet .
Portugal kan av sina finska föregångare lära sig hur det inte skall gå till .
Det är mycket viktigt att Europaparlamentet och kommissionen gör gemensam sak vid den här regeringskonferensen .
De har i många fall samma intressen och samma insikter .
En väsentlig del av den gemensamma insatsen måste i alla fall vara parlamentets medbeslutanderätt vid de kommande fördragsändringarna .
Av alla prioriteter så är det de som väger tyngst .
Vad anser kommissionen om det ?
Det betyder också att parlamentets ordförande och de två företrädarna måste kunna delta på en jämlik politisk nivå , alltså inte bara i arbetsgruppen utan på samma politiska nivå som kommissionen .
Det finns inget som helst skäl till att folkvalda företrädare skulle delta på en lägre nivå än kommissionen .
De grundliga reformerna är vi inte bara skyldiga de nya medlemsstaterna utan även oss själva .
Om vi låter Europa urvattnas på grund av utvidgningen så drunknar vi i vårt eget politiska träsk .
Herr talman !
Det finns dagar då jag verkligen inte förstår mig på detta parlament som finner en masochistisk njutning i självstympning .
Efter att på eget initiativ ha begränsat sitt deltagande i regeringskonferensen till två små platser avstår parlamentet i dag från att komplettera dagordningen för denna regeringskonferens .
Oavsett om det beror på svaghet eller dumhet , och ingen av dessa möjligheter är särskilt lysande det måste ni erkänna , överger vårt parlament , genom att skynda sig att yttra sig , den enda drivkraft som fördraget ger , dvs. att kräva en fullständig dagordning för regeringskonferensen innan man uttalar sig .
Varför skall vi brådskande rösta om detta yttrande i morgon den 3 februari när vi i vår styrkeposition kan vänta tills sammanträdet i Strasbourg öppnas den 14 februari , och på så sätt påtvinga rådet en dagordning som äntligen är fullständig och därmed enhetlig ?
Det krävs en hel del hyckleri för att dölja vår svaghet i dag .
Hyckleri för att i vår resolution allvarligt beklaga att regeringskonferensens dagordning inte är i nivå med vad som står på spel , medan vi med en skyldig naivitet gör allt för att undvika att tvinga fram denna ambitiösare dagordning .
Om det i slutet av denna regeringskonferens föreligger ett demokratiskt tomrum , då säger jag att de politiska grupper som velat ha denna brådska blir ansvarig för detta .
Vare sig man vill det eller ej kommer besluten att förskjutas mot de femton staterna i unionen , eftersom vårt parlament självt kommer att släcka den enda strålkastare som gjorde det möjligt att något lysa upp debatterna .
Jag uppmanar därför ledamöterna bland den enorma majoritet i parlamentet som i november ansåg att Europas framtid förtjänade bredare debatter än reliken från Amsterdam , att greppa sin vallfärdsstav och gå och övertyga sin regering om att vi måste utvidga denna regeringskonferens eftersom resolutionen från Europeiska rådet i Helsingfors tillåter det .
På grund av situationen i Österrike är denna dag en mörk dag för Europa .
Man inser då att demokratins seger aldrig är vunnen och att vi måste övertyga och övertyga igen .
För att bekräfta våra grundläggande värderingar är det brådskande att skriva dem och utöver denna regeringskonferens tror jag att vi är skyldiga Europa en konstitution .
Herr talman !
I det förslag till resolution som vi nu diskuterar krävs precis som tidigare att den kommande regeringskonferensen skall ha en bred dagordning med genomgripande reformer av institutionerna .
Som argument för detta används den kommande utvidgningen av unionen .
Jag är övertygad om att det är en felsyn .
Ett federalt och centralistiskt EU som styr alltmer i medlemsländerna har i själva verket sämre förutsättningar att utvidgas .
Ett flexibelt EU som koncentrerar sig på färre men viktiga områden och respekterar nationella olikheter och den nationella demokratin har bättre förutsättningar att omfatta betydligt fler länder .
I resolutionsförslagets punkt D krävs en mer samordnad och öppnare ekonomisk politik på EU-nivå .
Att tala om det är dock inte möjligt utan att samtidigt prata om den monetära unionen .
I den här texten sägs ingenting om de stora demokratiska och politiska problemen med valutaunionen och centralbanken - det är inte hållbart .
Vill man göra EU mer demokratiskt , måste EMU : s hela konstruktion omprövas .
Centralbanken måste ställas under politisk kontroll , så att valutapolitikens inriktning kan styras av politiska mål som hög sysselsättning och välfärd ; insynen i centralbanken måste förbättras för att detta skall bli möjligt .
Stabilitetspaktens stela och misslyckade monetarism måste omprövas och förkastas , för att vi skall kunna ha en enhetlig politik som sätter välfärdsmålen främst .
Fördragets artikel 56 , som förbjuder varje ingrepp i den fria rörligheten för kapitalet , valutaspekulationen , måste tas bort så att den skadliga valutaspekulationen kan hejdas genom politisk kontroll .
I flertalet EU-länder sitter i dag regeringar som domineras av socialdemokrater .
Det är anmärkningsvärt att ingen av dem kräver någon förändring i valutaunionens inriktning , nu när de har möjligheten .
Det skadar ju också trovärdigheten , när man påstår att valutaunionen skulle kunna utgöra en motvikt mot det globaliserade kapitalet .
I resolutionen kräver man att Europaparlamentet skall få ökat inflytande över regeringskonferensen .
Det är emellertid viktigt att understryka att regeringskonferensen är och skall vara en konferens mellan medlemsstaterna .
Det är medlemsländernas parlament , eller folk i folkomröstningar , som skall styra fördragets utveckling .
Det är därför uteslutet att Europaparlamentet ges något formellt inflytande i förhandlingsprocessen eller ratificeringen .
Herr talman !
Utskottet för konstitutionella frågor har föreslagit en text som i allt väsentligt är positiv , som jag kommer att rösta för , även om jag själv föreslog många ändringsförslag .
Det som under alla omständigheter har hänt under senare tid visar att alla de som riktade kritik mot hur utvidgningen och revideringen av fördragen planerades hade rätt .
Man kan inte utvidga unionen med 28 nya medlemmar utan att ta upp frågan om Europa har några principer , några gemensamma värderingar , om Europa reduceras till ett ekonomiskt frihandelsområde eller om det i stället har större ambitioner än så : att vilja vara en övernationell union , på ett sätt som måste definieras , som vill lägga ut ett nytt spår i världen mot humanitet och demokrati .
Det är detta vi önskar och menar när vi kräver en europeisk konstitution .
I stället har ändringen av fördragen begränsats till en revision av vissa interna regler , en nödvändig och viktig revision , men en som inte besvarar den grundläggande fråga som ställts : vad är Europa , vilka är dess gemensamma principer och därmed också dess mål och gränser ?
Men politiken hämnas och även om den kastats ut från fönstret i en debatt om en begränsad dagordning , så kommer den i själva verket tillbaka genom bakdörren , och i fallet Österrike genom ytterdörren , för i Österrike kommer ett parti till makten som tycks verka för intolerans , främlingsfientlighet , olika former av rasism .
Och det handlar inte om banden med det förflutna , detta är ett problem inför framtiden , och inget kunde vara felaktigare än att vi i den här frågan splittras mellan höger och vänster .
Jag tillhör en värld , de liberala katolikernas värld , som inte hör till vänstern men som står lika fast när det gäller försvaret av värden som tolerans , de gemensamma europeiska värderingarna , som alla andra och som vägrar ha något att göra med strömningar som förnekar sådana värden .
Rådet gjorde rätt som tog upp den här frågan i Europa och i världen och om vi inte fäster dessa värden i ett fördrag om grundläggande rättigheter , i en europeisk konstitution , så bygger vi upp ett Europa som inte har några fasta och hållbara grundvalar .
Jag vet , kommissionär Barnier - eller åtminstone så tror jag mig veta - att ni och samtliga företrädare för det portugisiska ordförandeskapet delar dessa värderingar : utnyttja de öppningar som kom från konferensen i december för att ta upp dessa frågor och dessa principer , för endast så kan vi konstruera ett hållbart Europa .
Herr talman !
Jag befinner mig i den glädjande situationen att jag kan hänvisa till ett par betydelsefulla inlägg från en liten grupp av nordiska skeptiker och motståndare till den våldsamma och övergripande integrationsprocess som i grunden hotar hela det demokratiska Europa .
Jag tänker på inläggen från Bonde och Sjöstedt , i vilka de påpekar att processen innehåller en rad förhållandevis aningslösa men tveklöst rationella och maktdikterade åtgärder i riktning mot ett centralistiskt och federalt EU .
De tog helt riktigt upp problemet med den monetära unionen och den centralistiska styrningen och ställde några alternativa demokratiska principer mot denna .
Jag kan tillfoga att all rationell politisk agitation i mitt hemland , Danmark , går ut på att när vi utvidgar kretsen av EU-länder till detta gigantiska antal , vi utvidgar alltså bredden , så kan vi inte samtidigt integrera mer på djupet - alltså genomföra en mer intensiv kvalitativ integration mot Europas förenade stater .
Men det är precis det som sker .
Vi har i samband med varje geografisk utvidgning av EU : s område sett att utvidgningar på bredden har följts upp av intensiva utvidgningar på djupet , och det är precis det som utskottets resolutionsförslag handlar om , särskilt punkt 7 i vilken det står att man skall ha en mer omfattande integration på djupet , och mot bakgrund av de senaste dagarnas utveckling kan man fråga sig vad vi egentligen skall ha dessa regeringskonferenser och fördragsändringar till , när regeringscheferna - i realiteten ministerrådet - fattar beslut i förhållande till en självständig medlemsstat , vilket innebär att man intervenerar i denna medlemsstats demokratiska process .
Man kan tycka vad man vill om Jörg Haider , och personligen tycker jag att han är en mycket farlig politisk person , men man kan ju inte intervenera i ett självständigt och vänligt sinnat lands demokratiska process .
När vi genomför regeringskonferenser och bedömer om vi skall genomföra fördragsändringar , måste vi ta hänsyn till att EU utvecklas varje dag , även i strid med fördraget som vi just har sett .
Jag hälsar kommissionär Barnier och det portugisiska ordförandeskapet välkomna här denna eftermiddag .
Den 14 februari inleds regeringskonferensen som skall avslutas i slutet av år 2000 .
Detta är en stor uppgift men den kan genomföras .
Jag tror att man allmänt inom alla grupper är överens om här denna eftermiddag att dagordningen i Helsingfors inte kommer att räcka till för att man skall hinna med det nödvändiga reformarbetet för att förbereda Europa inför utvidgningen .
Med andra ord vi måste täcka mer än vad som man har kallat de viktiga " Amsterdamresterna " .
Dessa innefattar utökad användning av omröstning med kvalificerad majoritet - i mitt land godkänner vi det , men inte när det gäller beskattningsfrågor - ny röstviktning i rådet för att gynna större stater samt antalet kommissionärer i ett utvidgat Europa .
Vad gäller den sista punkten vill Irland behålla rätten att nominera en fullvärdig och likvärdig ledamot av kommissionen utan hänsyn till det antal medlemsstater som ansluter sig .
Vi är beredda att överväga en ny röstviktning i ministerrådet , under förutsättning att de större medlemsstaterna är villiga att gå med på att varje medlemsstat får en fullvärdig och likvärdig ledamot i kommissionen .
Jag tror att jag talar för många mindre länder när jag hävdar den speciella åsikten .
Under regeringskonferensen behöver vi även debattera om en eventuell uppdelning av fördragen i två delar - en policydel och en konstitutionell del .
Vi kan godta uppdelningen av fördragen under förutsättning att det inte skulle begränsa den kontrollmöjlighet de mindre medlemsstaterna hade om omförhandlingen av fördragets alla politikområden .
Med andra ord om vi inte är helt företrädda i kommissionen kommer vi inte att kunna medverka i politiska diskussioner .
Således bevakar vi hela den frågan ytterst noga .
Vi ser fram emot stadgan om grundläggande fri- och rättigheter och att se dess innehåll .
I Amsterdamfördraget , herr talman , fastställs antalet ledamöter i Europaparlamentet till 700 och en debatt behövs i detta parlament om hur det antalet skall fördelas inom ett utvidgat Europa .
Herr talman !
Jag rekommenderar varmt att vi röstar igenom Dimitrakopoulos och Leinens resolution .
I resolutionen uttrycks tydligt såväl vår besvikelse över dagordningens otillräcklighet som vår vilja att regeringskonferensen skall klaras av så snabbt som möjligt .
Det framkommer för övrigt av den positiva tidtabell som vi har beslutat om .
Jag anser att Europaparlamentet , med de nuvarande fördragsreglerna , inte skulle ha mycket att vinna på en konfrontationspolitik .
Tvärtom bör vi koncentrera oss på att utarbeta övertygande förslag för de nödvändiga reformerna , i samarbete med kommissionen , vars förslag är värdefulla .
Vi måste utnyttja dialogen på alla politiska nivåer , inbegripet , naturligtvis , dialogen på de nationella parlamentens nivå .
Därigenom kommer vi att skapa ett samarbetsklimat som påverkar reformens kvalitet positivt .
Parlamentets företrädare på regeringskonferensen bör göra klart för förhandlingsparterna att vi framför oss , med de institutionella förändringarna för unionen , har ansvaret för unionens konstitutionella utveckling .
De måste därför inse att man inte beslutar om frågor av detta slag enbart med köpslagningslogik .
Frågorna för denna regeringskonferens är väldigt känsliga .
Det är möjligt att det är lätt för oss att lägga fram lösningar , frågan är dock hur bra dessa lösningar klarar av historiens granskning .
Jag vill betona två punkter som kan ge upphov till spänningar .
Den ena gäller den balans som fram till i dag har bevarats mellan de stora och de små staterna .
Europa är inte , och kan inte heller bli , en klassisk federal stat .
De lösningar som vi väljer måste ligga i linje med Europeiska unionens grundläggande logik , som är en förening av stater och den förening av folk .
Det andra området där det finns risk för kollisioner är svårare .
Vi kräver av den framtida europeiska unionen , på grund av den förestående ökningen av antalet medlemmar , att organen skall vara effektivare .
Det betyder att de skall fungera enklare och snabbare .
Europeiska unionen är dock av sin natur - och kommer så att förbli - en sammansatt och komplex flerstatlig institution .
Möjligheter till påskyndande och förenkling existerar .
Naturligtvis existerar de , men det finns gränser .
Om dessa gränser överskrids på grund av en ensidig effektivitet , kommer Europeiska unionens rättsliga grund att ha brutits ned .
Jag är emellertid optimistisk .
Herr talman !
Regeringskonferensens mandat måste utvidgas .
Den viktigaste frågan som bör läggas till är unionens interna differentiering .
Det är beklagligt att man knappt ens här i Europaparlamentet än så länge alls satt sig in i unionens interna differentiering som ändå är nödvändig för att unionen skall kunna utvidgas på det sätt som beslutats .
Kommissionens förre ordförande Jacques Delors har i offentlighetens ljus på nytt lyft fram tanken om en europeisk konfederation .
Han har också talat om att avant garde-länderna som ligger i täten för integrationen borde kunna gå framåt i snabbare takt än de andra och att de för klarhetens skull borde ha egna institutioner .
Kommissionens nuvarande ordförande Prodi och höge representanten Solana har framfört liknande tankar .
Europeiska liberala , demokratiska och reformistiska partiets grupp tog ställning till unionens interna differentiering genom en ståndpunkt som gruppen godkände i november i fjol och där man för Europeiska unionen föreslog ett system av cirklar med en gemensam medelpunkt , " en lökmodell " .
I nästa resolution om regeringskonferensen måste parlamentet på allvar sätta sig in i frågan om differentiering och flexibilitet .
Såväl utvidgningen som integrationens landvinningar är hotade om vi inte kan skapa ett system av cirklar med en gemensam medelpunkt .
Mina kollegor Frassoni och Onesta har redan ganska skeptiskt tala om några aspekter av den aktuella frågan .
Jag vill tillägga att jag är bekymrad över frågan om subsidiaritet , inte bara mellan union och medlemsstater utan mellan medlemsstater och deras egna internt självstyrande regioner .
Denna fråga har fått otillräcklig uppmärksamhet och här finns många bekymmersamma frågor .
Jag vill särskilt fästa er uppmärksamhet på en av utvidgningens följder för detta parlament .
Maximalt 700 har föreskrivits som den högsta antal som detta parlament kan bestå av utan risk och för att kunna förbli en rådgivande församling .
Om man tillämpar den nuvarande principen för avvikande proportionalitet , sex platser för varje stat och sedan en plats för varje halvmiljon innevånare har man redan situationen där Luxemburg med 367 000 innevånare har fler ledamöter i denna kammare än Wales som är en delvis självstyrande region i Förenade kungariket .
Skottland , med en befolkning på 5 miljoner , har åtta platser i denna kammare för ögonblicket ; Danmark och Finland , med samma befolkningssiffra , har sexton .
Vad kommer att hända om vi bibehåller en gräns vid 700 och för in 26 procent mer befolkning med tiden och sedan antar kommissionens som jag anser dåligt övertänkta förslag att det borde bli en europeisk kandidatlista .
Vad kommer att hända med ett land som Skottland , som jag företräder här ?
Det kommer att bli helt osynligt !
Ledamöter i denna kammare bör under dessa omständigheter inte alls bli överraskade om människor i Skottland och andra sådana länder vad gäller dessa diskussioner efterfrågar om utvidgning inte också borde innebära att nya medlemsstater inifrån redan existerande medlemsstater skall kunna ansluta sig .
En växande opinion i Skottland är av den åsikten .
Herr talman , herr rådsordförande , herr kommissionär !
Dagens debatt har en särskild politisk betydelse .
Det är inte fråga om att debattera innehållet , vare sig de punkter som redan finns med i dagordningen eller de som vi hade velat ha med , utan vi skall tala om vad Europaparlamentet anser om kallelsen till regeringskonferensen .
Och här finns inga nyheter , förutom en : att Europaparlamentet , i den här formen och genom sitt godkännande i morgon , valt en positiv strategi så att regeringskonferensen får en omfattande dagordning .
Genom sina ledamöter och talmannen visar man också sin vilja att bidra och berika en slutlig lösning av granskningen av fördraget .
Man ser positivt på kallelsen till regeringskonferensen , men är mera kritisk till dagordningens innehåll , vilket är helt naturligt .
Just nu är den institutionella ramen klar .
Det portugisiska ordförandeskapets positiva ståndpunkt och ambitioner är kända , Europaparlamentets ståndpunkt känner vi också till , kommissionen har just utarbetat ett dokument där man också klargör några av sina ståndpunkter , några anges som valmöjligheter , vilket gör att Europeiska rådet , om man använder sig av fotbollsjargong , " nu har bollen " .
Därför , herr talman och min käre vän Seixas da Costa , är min fråga följande : utan att vilja veta mera än det som vi just nu bör veta för att inte misskreditera det gemensamma målet så skulle jag , inom ramen för de resultat som uppnåtts efter den rundtur genom huvudstäderna som ni företagit och enligt er synpunkt , vilja veta om det finns några faktorer som kan bistå oss och vara oss till hjälp i vårt lobbying-arbete för bättre receptivitet och större inflytande över de nationella regeringar som är mest ovilliga att inkludera fler punkter på regeringskonferensens dagordning .
Min andra fråga riktar sig till kommissionär Barnier .
Den har att göra med kommissionens initiativ .
Jag var en av kritikerna : Jag tyckte att kommissionen borde ha gått längre vid Europeiska rådets möte i Helsingfors .
Jag tycker emellertid också att kommissionen har gjort ett utmärkt arbete , oberoende av om det överensstämmer eller inte med de lösningar som presenteras i det dokument som antogs den 26 .
Varför nöjer sig kommissionen med left overs från Amsterdam , eventuellt med en eller annan punkt till ?
Varför nöjer man sig med att nämna andra frågor som kan inkluderas , det vill säga dokumentet om de grundläggande rättigheterna eller frågor som berör den gemensamma utrikes- och säkerhetspolitiken ?
Därför vill jag uppmana kommissionen att , på samma sätt som när man på allvar tog tag i de förslag som vi redan känner till , gå händelserna i förväg och sätta igång och arbeta på de frågor som kanske längre fram kommer att ingå i dagordningen och därmed bidra till deras framgång .
Avslutningsvis , herr talman , vill jag lyckönska det portugisiska ordförandeskapet .
Uppgiften är inte lätt men jag vet att den är i goda händer .
Herr talman !
Påståendet att Europeiska unionen står i ett vägskäl innebär inget nytt .
Det är ett påstående som har upprepats vid flera tillfällen .
Men den här gången är det sant : vi har infört - något som är oerhört positivt - den gemensamma valutan och nu står vi inför en utvidgning .
Frågan är bara : skall vi vara förberedda eller ej när vi närmar oss en utvidgning ?
Är vi på väg att utvidga utan att gå grundligt tillväga eller är det just det vi gör genom att utvidga ?
Det är det som är frågan och dit leder varje diskussion beträffande regeringskonferensen , dess dagordning och metoder .
Det är uppenbart att rådet för ögonblicket inte har valt att utvidga genom att gå grundligt tillväga .
Det innebär en fara för utvidgningen .
Farligt , sett ur perspektivet av en politisk union , och givetvis svårt att förstå för allmänheten .
I rådet bör man vara medveten om att man måste gå betydligt längre på nästa regeringskonferens , om man i framtiden vill ha en väl förberedd utvidgning av Europeiska unionen .
Rådet rådfrågar oss och parlamentet lämnar sina synpunkter .
Vi vill ha en regeringskonferens , men inte denna .
Är det nödvändigt med en regeringskonferens ?
Ja , naturligtvis .
Men inte den här typen av regeringskonferens .
Man måste gå betydligt längre vad dagordningen beträffar , man måste vara betydligt djärvare i de frågor som tas upp under regeringskonferensen som måste erbjuda en ökad insyn och demokrati .
En ökad demokrati innebär att Europaparlamentet i högre grad tillåts medverka , att kommissionen i större - ja i större - utsträckning får utöva sin initiativförmåga .
Och givetvis att tydliga mål sätts upp .
Den funktionalistiska metoden har spelat ut sin roll , på gott och ont .
Så här långt har vi kommit med den funktionalistiska metoden .
Har vi uppnått några resultat ?
Jo då , men det gäller att ta ett kvalitativt språng , och det innebär i politiska termer , herr tjänstgörande rådsordförande , , att övertyga gemenskapens medlemmar om att det värsta vi nu kan göra är att inte uppnå målet .
Herr talman , mina damer och herrar parlamentsledamöter !
På det här stadiet och efter den debatt som jag lyssnat till mycket uppmärksamt och med stort intresse , skulle jag vilja göra några kommentarer som kompletterar de riktlinjer eller anföranden som jag redan haft äran att hålla för er de senaste veckorna , vid ordförande Prodis sida .
Herr talman , mina damer och herrar !
Era två föredragande , Dimitrakopoulos och Leinen , föreslog i det betänkande de lagt fram efter ett mycket exakt och seriöst arbete , att parlamentet skulle anta ett formellt yttrande enligt artikel 48 i fördraget och att regeringskonferensen med hjälp av detta yttrande effektivt kan inledas den 14 februari , såsom det portugisiska ordförandeskapet föreslagit .
I vårt ställe , och efter att utifrån samma artikel 48 i fördraget ha åstadkommit det yttrande som förväntades från kommissionen , är vi glada över att konferensen därför kan inledas , för övrigt tidigare än vad man ursprungligen tänkt .
Vi vet , jag vet , att alla de veckor vi har framför oss kommer att vara nyttiga veckor .
Jag skulle bara vilja göra några kommentarer efter att ha läst detta förslag till yttrande , och efter att ha lyssnat till talarna från de olika grupperna .
Mina damer och herrar !
Till att börja med förstår kommissionen den oro som flera av er uttryckt när det gäller omfattningen dagordningen för konferensen .
Jag förstår denna oro , denna fruktan att dagordningen skall vara alltför tvingande och det förefaller mig ändå som om vi kan arbeta , såsom jag sade till utskottet för konstitutionella frågor efter Helsingfors , på grundval av detta mandat från Helsingfors .
Det är just i den andan och inom ramen för detta mandat , men genom att använda alla fraser , allt som står skrivet mellan raderna i detta mandat , som kommissionen själv arbetat för sitt eget yttrande .
Vi är inte begränsade till vad man , för övrigt oriktigt , kallar de tre resterna .
Precis som Richard Corbett tycker jag inte heller om ordet " rester " , som ger en känsla av att det handlar om tre små frågor eller frågor utan betydelse .
Det handlar om tre mycket allvarliga , viktiga och svåra frågor , så svåra att det kollektiva politiska modet svek oss för att behandla dem på djupet i Amsterdam .
När det gäller oss - jag svarar Seguro , som nyss oroade sig på den punkten - har vi inte nöjt oss med dessa tre frågor , även om jag anser att de är de viktigaste och att vi nu måste behandla dem .
De är de första , de är inte de enda frågorna , herr parlamentsledamot , som konferensen måste behandla .
Vi har behandlat andra frågor och vi har tagit upp idén att andra frågor borde behandlas under denna konferens , om det portugisiska ordförandeskapet till att börja med vill , och sedan det franska , med tanke på allvaret i det vi upplever före utvidgningen .
Vi är beredda att göra det , vare sig det handlar om stadgan om de grundläggande rättigheterna , där arbetet påbörjats , eller om GUSP och de institutionella konsekvenserna av förhandlingarna som ägt rum om försvarspolitiken , eller om en mycket svår fråga som vi fortsätter att arbeta med , nämligen omorganisationen av fördragen .
Jag har hört många kommentarer om kommissionens yttrande , som tog upp alla dessa frågor och som behandlade många av dem grundligt , inbegripet exakta demonstrationer av förslag till nya artiklar , men ingen har sagt att vi befinner oss utanför mandaten från Helsingfors .
Det är därför beviset på att man samtidigt som man respekterar mandatet kan , genom att använda allt det som skrivits i mandatet och alla de öppningar det innehåller , gå till botten med frågorna .
När det gäller Europaparlamentets deltagande i arbetet med konferensen tror jag att minister Seixas da Costa är överens med mig , eftersom vi har en gemensam erfarenhet , när jag säger att det skulle vara fel av er att strunta i nivån med diskussions- och förhandlingsgruppen där era två företrädare , professor Tsatsos och Elmar Brok , kommer att arbeta .
De sista skiljeförfarandena kommer naturligtvis , såsom alltid är fallet i varje institutionell förhandling , att äga rum och jag tror att det är bra , inom rådet och framför allt bland stats- och regeringscheferna , som kommer att ha framgången för denna konferens i sina händer .
Jag vill också i förbigående påpeka att kommissionens ordförande Prodi ingår i rådet och han har för avsikt att utnyttja denna plats och denna roll , vid stats- och regeringschefernas sida , bl.a. under slutperioden .
Men vi måste noga förbereda detta arbete i rådet .
Mina damer och herrar parlamentsledamöter !
Vi får alltså inte bortse från detta förberedelse- och förfiningsarbete som jag , genom min erfarenhet från Amsterdam , vet är mycket viktigt och användbart , och man skall inte bara nöja sig med tekniska preciseringar .
Jag tror att de personliga företrädarna för utrikesministrarna , era två företrädare och jag själv som företrädare för kommissionen , kommer att gå till botten med saken , men det blir senare , på en annan nivå , där vi också skall delta , som de sista skiljedomarna kommer att genomföras .
Under hela denna konferens , mina damer och herrar , är det inte bara ställningen för förhandlarna som är viktig , utan kvaliteten i vad de säger .
Och jag vill än en gång med tanke på mina erfarenheter från Amsterdam inför parlamentet upprepa , oavsett vilken tvetydig eller svag ställning de två företrädarna från Europaparlamentet har , att före Amsterdam var kvaliteten i vad Guigou och Brok sade av stor betydelse i denna förhandling .
Jag är säker på att det blir samma sak när det gäller mig , på min plats , och jag skall se till att idéerna från era två företrädare uppmärksammas och respekteras under hela förhandlingen .
Jag är säker på att Europaparlamentet då inte blir åskådare till denna förhandling , på samma sätt som kommissionen inte heller blir det .
Mina damer och herrar parlamentsledamöter !
Vi väntar därför med stort intresse på ert yttrande senare där ni kommer att precisera prioriteringar och konkreta förslag från parlamentet inför förhandlingen .
Det är av stor vikt att de två europeiska institutioner som kommer att närvara vid dessa förhandlingar , kommissionen respektive Europaparlamentet , vid sidan av rådets medlemmar , alltid och varje dag tydligt förklarar för medborgarna i unionen vilka frågor som står på spel under denna konferens och vilka svar vi förespråkar som europeiska institutioner , med ansvar för att se till att denna utvidgade union fungerar korrekt och i allas intresse .
Mina damer och herrar parlamentsledamöter !
Under de kommande månaderna kommer alltså kommissionen att arbeta i nära samråd , och på ett intelligent sätt , med era två företrädare , professor Tsatsos och Elmar Brok , för att närma våra ståndpunkter till varandra , om det behövs .
Sannolikt kommer våra ståndpunkter och våra positioner inte alltid att vara desamma , det kommer säkerligen att föreligga skillnader , vilket är normalt .
Det som är viktigt , är att det föreligger enhetlighet , det är för att arbeta med denna enhetlighet som jag redan från början engagerat mig i mitt ämbete inom kollegiet .
Vi har alltså strävan och ambitionen , i ett mycket stort antal frågor , att befinna oss på samma våglängd och höja förhandlingen .
Det är ingen tillfällighet eftersom , jag upprepar det , det förefaller som om vi har samma ambition för denna förhandling och vi känner tillsammans att den verkligen utgör en sanningens minut för Europeiska unionen .
Herr ordförande !
Jag skulle slutligen litet snabbt vilja göra tre kompletterande kommentarer .
Till att börja med för att lyckönska och tacka ordförande Napolitano och utskottet för konstitutionella frågor för det mycket starka och originella initiativ som togs i går genom att samla kvalificerade företrädare från de nationella parlamenten , utskottet för konstitutionella frågor och kommissionen för en första gemensam debatt .
Denna dialog mellan de nationella parlamenten , Europaparlamentet och oss själva är mycket viktig .
Jag sade för övrigt att jag skulle ta mitt ansvar genom att själv besöka samtliga nationella parlament .
I morgon kommer jag att vara i London .
Om två veckor är jag i Berlin .
Om tre veckor i Paris , och sedan skall jag fortsätta , huvudstad för huvudstad , att i min tur delta i denna dialog .
Jag finner det mycket positivt och jag ville tacka er för att ni tagit detta initiativ .
Ytterligare några ord för att tacka det portugisiska ordförandeskapet och särskilt herr Seixas da Costa , för hans voluntarism .
Det han nyss sade visar tydligt på den voluntarism och den oro som också han har : det portugisiska ordförandeskapet kan inte vara ett mellanliggande ordförandeskap .
Det är detta ordförandeskap som skall inleda förhandlingen .
Vi vet mycket väl att den inte kan avslutas under dessa sex månader och att det franska ordförandeskapet sedan skall ta över , med förhoppningen att det skall avsluta förhandlingen innan år 2000 är slut .
Och inte bara avsluta , utan också lyckas med den , vilket inte är riktigt samma sak .
Att avsluta en förhandling är inte detsamma som att lyckas med den .
Ordförandeskapet kommer att ha överlämnats , men under vilka förhållanden detta överlämnande sker av er själv , herr ordförande , och av det portugisiska ordförandeskapet , blir mycket viktigt , liksom hur det sker .
Det är det arbete som vi skall genomföra tillsammans , och bl.a. med impulser från er , under några månader , vilket är mycket viktigt .
Vi hyser stort förtroende för er och vi har stora förväntningar på det sätt som det portugisiska ordförandeskapet , från ett litet land - men även om man är liten kan och bör man ha stora ambitioner - kommer att genomföra denna uppgift .
Efter att ha lyssnat till premiärminister Guterrez , utrikesministern och er själv , hyser jag detta förtroende för ambitionen hos det portugisiska ordförandeskapet och det mycket voluntaristiska sätt som det kommer att föra denna förhandling på .
Ordförandeskapet kan under dessa månader räkna med kommissionens partnerskap .
Slutligen , jag upprepar det , har vi en mycket stor ansträngning framför oss för att popularisera frågorna i denna förhandling .
Det är svåra frågor .
Det är frågor om institutionell politik och mekanik som inte alltid är lätta att förklara .
Det är ytterligare en anledning till att ledamöterna i Europaparlamentet , ministrar och kommissionärer bör ägna litet tid åt att förklara för medborgarna och bedriva en offentlig debatt .
Kommissionen kommer för sin del att ta initiativ , mina damer och herrar , till att inleda och föra denna debatt .
 
Utförande av tjänster över gränserna Nästa punkt på föredragningslistan är gemensam debatt om följande betänkanden : A5-0007 / 2000 av Berger för utskottet för rättsliga frågor och inre marknaden om förslaget till Europaparlamentet och rådets direktiv om utstationering av arbetstagare från tredje land i samband med tillhandahållande av tjänster över gränserna .
( KOM ( 1999 ) 3 - C4-0095 / 1999 - 1999 / 0012 ( COD ) ) A5-0012 / 2000 av Berger för utskottet för rättsliga frågor och inre marknaden om förslaget till rådets direktiv om en utvidgning av friheten att tillhandahålla tjänster över gränserna till att även omfatta tredjelandsmedborgare som har etablerat sig inom gemenskapen ( KOM ( 1999 ) 3 - C4-0096 / 1999 - 1999 / 0013 ( CNS ) ) .
Herr ordförande , herr kommissionär , värderade kolleger !
Till att börja med måste jag be om ursäkt för att jag är litet hes i dag , men som österrikisk ledamot har man haft mycket att förklara och tala om i dag .
Jag vill först tacka kommissionen så hjärtligt för det initiativ som den har tagit , och för de båda förslag till direktiv som vi diskuterar här i dag .
Den åtgärdar därmed två graverande brister på den inre marknaden som är av stor betydelse för det europeiska näringslivet och för 5 miljoner tredjelandsmedborgare i Europeiska unionen , vilka är här som arbetstagare eller som individer .
Dagens situation , och det bör man än en gång betänka , ser ut så att det i fråga om arbetstagarna visserligen föreligger domar från EG-domstolen , i synnerhet domen som gäller Rush Portuguesa och van der Elst .
De har visserligen klarlagt att friheten att tillhandahålla tjänster måste medge att man använder sig av tredjelandsmedborgare som arbetstagare för gränsöverskridande tjänster , och detta även utan att kunna utverka arbetstillstånd .
Frågan om viserings- och uppehållsvillkor fördes inte utförligen på tal , och inte heller medlemsstaterna kunde sedan förklara denna fråga .
Men inte heller med hänsyn till bortfallet av arbetstillståndet har alla medlemsstater hållit sig till domstolens domslut utan upprätthåller fortfarande i dag en mängd otillåtna barriärer för gränsöverskridande tjänster , barriärer som ofta är omöjliga att övervinna , i synnerhet för små företag .
För de egna företagarna ser situationen så ut att gemenskapens nuvarande regelverk inte föreskriver någon rätt för tredjelandsmedborgare att utföra gränsöverskridande tjänster .
Här behöver man i varje fall en rättsakt .
Båda förslagen till direktiv syftar till att underlätta friheten att tillhandahålla tjänster för EU-företag .
Det handlar inte om nya rättigheter för tredjelandsmedborgare , som efterbildar den fria rörligheten .
Alla bestämmelser , inresa och frågor som gäller uppehållet , skall betraktas som tillägg till denna frihet att tillhandahålla tjänster .
Tillsammans med utskottet för rättsliga frågor och den inre marknaden anser jag därför att den av kommissionen valda rättsliga grunden är riktig och att den motsatta åsikt som företräds i utlåtandet från rådets rättstjänst inte är tillämplig .
Jag ser därför inte heller något verkligt hinder för att båda förslagen till direktiv snabbt skall kunna vidarebehandlas i rådet .
Jag tror också att de av parlamentet föreslagna ändringarna bör göra att direktiven lättare blir antagna i rådet , jämfört med kommissionens förslag .
Många av våra ändringar går tillbaka till betänkligheter som även yttrats i rådet , och vi försöker att förena dessa betänkligheter med det uppdrag som gällande rätt och ekonomiskt förnuft ger oss .
Även med tanke på acceptansen i rådet kan jag bara vädja till kommissionen att så snart som möjligt fullständigt överta de ändringar som parlamentet antagit , även om de delvis avviker avsevärt från kommissionens ursprungliga förslag .
Jag är fast övertygad om att vi på denna grundval lättare kan uppnå enighet i rådet .
Nu till de viktigaste ändringarna som vi föreslår .
En väsentlig skillnad består i att vi i stället för ett system med frihet att tillhandahålla tjänster plus anmälning av varje enskilt uppdrag inte längre räknar med möjligheten att man för varje enskilt uppdrag skall kunna begära att det i förväg anmäls till det mottagande landet .
Detta system förefaller oss oanvändbart i praktiken .
Som kompensation för detta måste dock , innan EG-kortet för tillhandahållande av tjänster ställs ut , alla eventuella hinder ha undanröjts , och gentemot kommissionens förslag måste skärpta villkor ha uppfyllts för att EG-kortet för att tillhandahålla tjänster skall kunna ställas ut .
Kraven på vederbörlig sysselsättning , legalt uppehåll och försäkringsskydd måste finnas inte bara vid tidpunkten då EG-kortet ställs ut , utan under hela kortets giltighetstid , plus tre månader därefter .
Därigenom bör den mottagande staten ha en garanti för att arbetstagaren respektive den egna företagaren efter fullgjort uppdrag också återvänder till den stat han kommer från , och i händelse av sjukdom och olycksfall täcks av försäkringar .
Inresan och situationen som rör uppehållstillståndet skall också ha klarlagts innan kortet för tillhandahållande av tjänster ställs ut , nämligen inom ramen för ett överklagandeförfarande .
Vi föreskriver att EG-kortet för tillhandahållande av tjänster inte måste begäras för alla medlemsstater , utan att det också kan begäras för enskilda medlemsstater .
Jag tror att detta system också bättre motsvarar de praktiska behoven .
Samma sak hoppas jag man åstadkommer genom förslaget att sänka minimilängden för den tidigare sysselsättningen till tre månader , och att inrikta giltighetstiden för kortet för tillhandahållande av tjänster beroende på längden på den tidigare sysselsättningen på ett flexibelt sätt .
Men vi anser fortfarande att den maximala giltigheten för kortet för tillhandahållande av tjänster skall ligga vid 12 månader .
Vad gäller de egna företagarna föreslår vi också , som tillägg till de redan beskrivna ändringarna , att etableringskriteriet måste skärpas och att vi föreskriver en möjlighet att bemöta ett eventuellt missbruk på grund av falskt egenföretagande .
Jag vill också kort gå in på föreliggande ändringsförslag , som går utöver ändringsförslagen från utskottet för rättsliga frågor och den inre marknaden .
Jag vill naturligtvis också säga att jag även i fortsättningen stöder de av detta utskott framlagda ändringarna , som antogs enhälligt i utskottet .
Jag har själv för min grupp lämnat in fyra ändringsförslag , som väsentligen hänför sig till det korrekta sättet att citera ett beslut från rådet .
Jag måste säga att jag här från parlamentets tjänsteenheter har fått ytterst motsägande uppgifter om hur nu detta beslut från rådet skall citeras korrekt ; endast med nummer , endast med datum , med båda , hur utförligt det skall citeras från rådets beslut .
Två ändringsförslag togs bort av tjänsteenheterna , eftersom man enligt uppgift redan tagit hänsyn till innehållit i dem i betänkandet .
Jag drar tillbaka de två ytterligare ändringsförslagen - det är ändringsförslag 18 i betänkandet om egenföretagarna och 21 om de anställda .
Jag kan bara vädja till talmanskonferensen att så snart som möjligt enas om hur man i fråga om kommittésystemet skall agera korrekt när det gäller citat .
Det skulle underlätta livet för föredragandena i denna kammare väsentligt i framtiden .
Det föreligger också ett ändringsförslag till båda betänkandena från kollegan De Palacio .
Jag måste tyvärr säga att jag inte kan stödja detta ändringsförslag , eftersom det skulle förändra substansen i de resultat som vi enhälligt uppnådde i utskottet för rättsliga frågor och den inre marknaden , och jag vill bibehålla det som vi i detta utskott efter långa diskussioner gemensamt kom fram till .
Avslutningsvis vill jag tacka alla kolleger som har bistått mig i utskottet för rättsliga frågor och den inre marknaden i dessa inte direkt lätta betänkanden .
I synnerhet vill jag nämna kollegan Wieland , som har den otacksamma rollen som medföredragande och långt utöver det vanliga tagit del i utformningen av detta betänkande med mycket bra och konstruktiva idéer , utan att få någon del av föredragandens lagerkrans .
Därför vill jag här särskilt nämna det ! .
( NL ) Herr talman !
Jag är glad att jag får tillfälle att efter anförandet av föredraganden , Berger , göra några inledande kommentarer varefter jag naturligtvis med allt det intresse som krävs skall lyssna till de följande talarna .
Om ni tillåter , herr talman , skulle jag sedan i slutet av debatten vilja ta upp de olika ändringsförslagen mer ingående .
Jag vill tala om att kommissionen gläder sig åt Europaparlamentets stöd för de två förslag för tillhandahållande av tjänster och arbetstagare från tredje land , vilka debatten nu gäller .
Jag är särskilt tacksam för det arbete som Berger lagt ner vid behandlingen av de här förslagen som ju är politiskt känsliga och som är en politisk utmaning .
Jag vill också tacka Palacio så mycket för hennes mycket viktiga bidrag som ordförande för utskottet för rättsliga frågor och den inre marknaden .
Kommissionen gläder sig särskilt åt parlamentets förslag om ett effektivare förfarande för utfärdande av kortet för tillhandahållande av tjänster .
När det finns möjlighet att ansöka om ett sådant kort för en eller flera eller för alla medlemsstater så blir förfarandet ännu flexiblare .
Kommissionen går också med på den föreslagna giltighetstiden för kortet .
Jag anser emellertid att en arbetsperiod på tre månader inte räcker som bevis för att en arbetstagare är etablerad i en medlemsstat .
Kommissionen kan också gå med på en bestämmelse för de fall då arbetskontraktet mellan tjänsteleverantören och arbetstagaren plötsligt upphävs .
Ett effektivt förfarande för utfärdande av kortet innebär att företag som tillhandahåller gränsöverskridande tjänster också verkligen kan utöva sina rättigheter på grund av den inre marknaden .
Vi tycker att det verkar överdrivet om andra medlemsstater får möjlighet att för utfärdandet av ett kort genomföra systematiska kontroller med avseende på den allmänna ordningen .
En medborgare från ett tredje land med en legal ställning måste ju också få komma in i andra medlemsstater .
Det hindrar inte dessa medlemsstater från att inom ramen för den föreslagna meddelandeskyldigheten vidta åtgärder med avseende på den allmänna ordningen .
Förslaget om att uppehållstillståndet i en medlemsstat borde vara tre månader efter kortets giltighetstid kan kommissionen inte heller godta .
Det är inte godtagbart att den berörda medborgaren från ett tredje land stannar längre i medlemsstaten efter det att tjänsterna tillhandahållits .
Därför stöder kommissionen i båda fallen ändringsförslag 22 av Palacio .
När det gäller det andra förslaget så inser kommissionen att det måste vara tydligt vad som menas med en egenföretagare och skall därför komma med en lösning i det ändrade förslaget .
Det var några inledande kommentarer om de viktigaste ändringsförslagen .
Jag hoppas att jag i slutet av den här debatten , när alla talare sagt sitt , får ytterligare tillfälle att ta upp de olika ändringsförslagen .
Herr talman , mina damer och herrar !
PPE-gruppen kommer med stor majoritet att rösta för ändringsförslagen från utskottet för rättsliga frågor och den inre marknaden och även den ändrade versionen under morgondagen .
Jag vill i mina utlägg inskränka mig till två betänkanden .
Det ena gäller frågan om vad detta direktiv över huvud taget skall verka för - verka för i dess egentliga betydelse .
Vi har för det första näringslivets och även de enskildas intressen .
I mina inlägg utgår jag till att börja med från att det handlar om en rättskaffens och rejält arbetande enskild .
För det andra har vi medlemsstaternas intressen , som med tanke på dem som berörs kanske också måste utgå från att det föreligger ett worst case .
Om vi tänker på den ena ytterligheten , medlemsstaternas intressen , så finns det säkert goda anledningar att sätta hindren för detta EG-kort relativt högt .
Sedan finns det anledning att trots detta EG-kort på ett tidigt stadium införa anmälningsplikt .
Om jag tänker på den andra ytterligheten , alltså så få hinder som möjligt , då riskerar jag att jag i fråga om detta förfarande över huvud taget inte kommer att få uppleva någon lagstiftning , eftersom medlemsstaterna då inte kommer att godkänna direktivet .
Resultatet blir alltså antingen att jag visserligen har ett direktiv för EG-kortet för tillhandahållande av tjänster , men , eftersom hindren för näringslivet är mycket höga , i själva verket inte har något EG-kort för någon .
I det andra fallet har jag inte alls något direktiv .
Ingetdera resultatet är tillfredsställande .
Kanske är detta också anledningen till , som man hör sägas , att förhandlingarna har hakat upp sig även i rådet .
Nu har vi försökt att åstadkomma ett mellanting mellan det ena intresset - ordre public - och det andra intresset , och att finna en så lätt lösning som möjligt .
Vi vill ha en lösning där vissa hinder för näringslivet byggs upp , men där man sedan , när dessa hinder övervunnits , uppnår en så smidig hantering som möjligt .
Vi vill därför att EG-kortet för tillhandahållande av tjänster begärs för en eller flera medlemsstater .
Om ett företag i Frankrike säger att man har en medarbetare som ständigt måste arbeta i Danmark och bara i Danmark , då skall detta EG-kort för tillhandahållande av tjänster också bara begäras för Danmark .
Då kommer de byråkratiska hindren för detta att vara lägre .
Som en motåtgärd vill vi dock att det inte längre skall finnas några fler tidiga anmälningsplikter , utan att arbetstagaren enbart skall ha med sig anledningen till arbetena i den andra medlemsstaten , till exempel i form av det avtal som ligger till grund för dem .
Därför måste jag också säga att jag till slut uttalar mig för ändringsförslagen från utskottet för rättsliga frågor .
Kanske finns det också hos kommissionen fortfarande kvar en viss rest av missuppfattning .
Vi vill att man uppnår en helt flexibel lösning .
Om en medlemsstat förklarar att man plötsligt har problem , eftersom personen har begått en stöld , man har problem , och detta EG-kort för tillhandahållande av tjänster är utställt för ens land , då kan det enskilda landet av de anledningar som finns i detta direktiv i viss mån dra tillbaka giltigheten för EG-kort , på ett flexibelt och intelligent sätt .
Låt mig också helt kort gå in på en annan sak .
De flesta som hittills befattat sig med direktivet är jurister .
Vi vet alla att det fortfarande finns olika beståndsdelar i fördraget , delvis mycket gamla beståndsdelar i fördraget , som fortfarande heter EG .
Vi vet att detta direktiv baserar sig på EG-rätt och inte på EU-rätt .
Men före valet verkade vi - rådet , kommissionen , parlamentet , pressen , fackföreningarna , organisationerna - för att detta Europa skall bli mer förståeligt för medborgaren .
Vi har ansträngt medborgarna genom att ändra EEG till EG till EU .
Nu har man förstått EU .
Vi gör oss själva och medborgaren en otjänst om vi nu döper den produkt som vi ger ut till EG-kort för tillhandahållande av tjänster och inte till EU-kort för tillhandahållande av tjänster .
För medborgaren är EU-världen intressant , det är den som gäller för honom .
Jag ber rådet och kommissionen att gå i den riktningen .
Herr talman !
Det har blivit senare än någon av oss trodde det skulle bli när vi planerade denna session så jag skall verkligen fatta mig kort .
En av orsakerna till varför vi är försenade är för att vi använde tiden tidigare i dag till att rätteligen framföra det fast förankrade motståndet i detta parlament mot varje form av främlingsfientlighet och rasism .
Detta direktiv handlar naturligtvis inte i sig självt direkt om det .
Det handlar om att se till den inre marknadens behov , att skapa flexibilitet och att agera på ett förnuftigt och flexibelt sätt för att skapa sysselsättning för människor från tredje land både som anställda och som egenföretagare .
Det handlar i sig själv också om att undvika att vara obefogat restriktiv mot främlingar bara för att han eller hon är en främling .
Vi välkomnar det och då vi anser att det är en förnuftig och riktig bestämmelse kommer vi att stödja den mest generösa versionen som vi anser är i överensstämmelse med lagstiftningen . .
( ES ) - Herr talman , herr kommissionär !
Jag vill börja med att poängtera det utmärkta arbete som Berger har gjort och även rent allmänt utskottet för rättsliga frågor och den inre marknaden , som har infört nyskapande idéer i detta direktiv som jag hoppas kommer att godkännas av kommissionen och rådet .
Jag har emellertid lagt fram ett ändringsförslag .
Fru Berger , i ert ändringsförslag 2 , skäl 6 , tar ni upp rättssäkerheten .
Den första punkt där vi har en avvikande mening är uppehållstillståndets förlängning med tre månader , för det skapar endast rättsosäkerhet .
Ni har - av naturliga skäl - uttryckt er oro , som bekräftats av Wieland , för möjligheten att en arbetstagare försvinner när dennes arbetstillstånd har löpt ut , men jag anser att ni samtidigt underlättar denna möjlighet i och med förlängningen med tre månader .
Om giltigheten för EG-kortet för tillhandahållande av tjänster upphör ett visst datum , bör den också upphöra det datumet .
Det är en förutsättning för rättssäkerheten .
Å andra sidan , vad beträffar punkt d ) i ändringsförslag 10 som åsyftar det första direktivet , nämner ni att en medlemsstat på grund av allmänhetens säkerhet eller bestämmelser om den allmänna ordningen , kan vägra erkänna kortets giltighet .
Redan nu sker kontroller som ex ante fastställs i artikel 4 i direktivet .
Det saknar betydelse för en arbetstagare inom Schengenområdet , för denne har redan genomgått en kontroll för att få resa in i den första medlemsstaten , och den andra medlemsstaten kan ex ante , om vissa skäl föreligger , neka denna arbetstagare inresa i landet .
Det finns därför ingen anledning att bevara denna rättsosäkerhet .
Om det inte rör sig om en Schengenstat så förutses den möjligheten i sista stycket i mitt ändringsförslag 22 , i alla avseenden och med det jag anser vara en bättre rättssäkerhet .
Staternas fria val som ni föreslår i punkt e ) i ert ändringsförslag 10 rimmar inte med texten i övrigt i ert utmärkta betänkande .
Därför uppmanar jag er kolleger att ta del av mitt ändringsförslag , och hoppas att vi i morgon kan komma fram till en lösning .
Av allt att döma tycks dessa två förslag införa vissa ändringar i förfarandena för att underlätta fri rörlighet i hela Europa och för att låta de nya domstolsfall som Berger refererade till i sitt öppningsanförande få effekt .
I fråga om Förenade kungariket tror vi emellertid att man där går längre än så på ett sätt som är oacceptabelt .
Delvis finns verklig substans delvis är det med hänsyn till den rättsliga grunden vad gäller Förenade kungarikets särskilda ställning .
Enligt de protokoll som finns i fördragen behåller Förenade kungariket sin egen gränskontroll .
Enligt det system som föreslagits på dessa lagstiftningsområden kommer medborgare i tredje land som vill flytta till Förenade kungariket att enligt de beskrivna förfarandena kunna göra detta med hjälp av ett servicekort utfärdat av en annan medlemsstat och därigenom kringgå landets gränskontroller .
Om det nuvarande gränskontrollsystemet i Förenade kungariket skall ändras bör den ändringen göras av Förenade kungarikets regering och parlament och inte i förbifarten genom det europeiska lagstiftningsförfarandet .
Av det skälet skall vi rösta mot båda dessa förslag .
Herr ordförande , herr kommissionär , mina damer och herrar !
Först vill jag tacka föredraganden och kollegan Wieland så hjärtligt för deras ansträngningar att så homogent sammanfatta de olika ändringsförslagen och de olika intressena i detta betänkande .
Dessa båda förslag bidrar till att genomföra en av de fyra kärnprinciperna för den inre marknaden , fri rörlighet för tjänster .
De nya bestämmelserna för gränsöverskridande tjänster kommer utan tvivel att förbättra både den inre marknadens funktion och företagens konkurrens- och handlingskraft .
De strikta ramvillkoren för utställandet av - och här citerar jag kollegan Wieland - EU-kortet för tillhandahållande av tjänster är oundgängliga , eftersom de tjänar till att förhindra missbruk , exempelvis illegal invandring och falska kontrakt .
Varför anser jag att direktivet är så nödvändigt ?
Av tre anledningar : På grund av den ekonomiska betydelse som arbetskraften från tredje land har i EU , på grund av företagens konkurrenskraft och på grund av den inre marknadens friktionsfria funktion .
Därför välkomnar jag å ena sidan den strikta ramen , och vädjar å andra sidan om att de lämpliga kontrollerna som medlemsstaterna genomför blir så effektiva och enkla som möjligt .
Min sista fråga , eftersom man alltid frågar mig om det , går till kommissionen : Kommer direktivet att bli prejudicerande för anslutningsförhandlingarna ?
Hur kommer artikel 1 ur er synpunkt att tolkas , eftersom detta spelar en viktig roll i anslutningsförhandlingarna och just för vårt land som gränsar till många nya länder ?
Herr talman , herr kommissionär , kolleger !
De företagare som hittills tvingades konstatera att två av de viktiga friheterna , nämligen fri rörlighet för personer och tjänster , inte gällde för dem var dock tvungna att gå igenom en oändlig byråkratisk immigrationsprocess i medlemsstater där en tjänst skulle tillhandahållas .
Det finns cirka tretton miljoner medborgare från tredje land som uppehåller sig i Europa .
Jag utgår från att , även om det inte är känt exakt hur många av dem som är företagare , deras antal säkert inte är litet .
Hittills har deras tillträde till hela Europeiska unionen inte reglerats genom gemenskapsrätten .
Syftet med de två aktuella förlagen till direktiv är att främja den fria rörligheten för tjänster på den inre marknaden genom införande av EU-kortet för tillhandahållande av tjänster .
Jag tycker det är viktigt att i det sammanhanget understryka att utfärdandet av ett sådant kort skall ske på ett flexibelt sätt , nämligen inom fem dagar efter att en enkel förklaring lämnats till den medlemsstat där tjänsten skall tillhandahållas och att , för att undvika missbruk , den här handlingen skall ha en begränsad giltighet och inte automatiskt kunna förlängas .
Jag har också med intresse tagit del av de invändningar som kommissionären fört fram här .
Efter att ha studerat de inlämnade ändringsförslagen har jag också konstaterat att vi i stor utsträckning kan godta dessa invändningar och därför skall anpassa hur vi röstar efter detta vid omröstningen i morgon .
Avslutningsvis skulle jag vilja tacka föredraganden Berger för den noggrannhet med vilken hon undersökt de olika ändringsförslagen och på det sättet givit sitt betänkande ett viktigt innehåll .
Jag tror att vi med det här betänkandet tagit ett nytt steg mot förverkligandet av den inre marknaden . .
( NL ) Herr talman !
Tack för att jag nu får tillfälle att mer specifikt gå in på de olika ändringsförslagen och i det sammanhanget skulle jag också vilja säga något till Lord Inglewood om den anmärkning han nyss gjorde .
När det gäller det första förslaget om arbetstagare från tredje länder så är kommissionen beredd att anta ändringsförslagen 2 , 11 , 12 , 15 , 16 och 22 .
Även ändringsförslagen 7 och 8 är godtagbara om utstationeringssituationen i ursprungslandet kan fastställas .
Kommissionen godtar också ändringsförslag 11 , förutom med avseende på den föreslagna perioden för tidigare anställning på endast tre månader .
Det har jag redan förklarat tidigare .
Även ändringsförslag 13 är välkommet om det härigenom införs ett flexibelt tillämpningsområde för kortet från en medlemsstat till alla medlemsstater .
Vad kommittésystemet beträffar så kan ändringsförslagen 14 och 21 också delvis godtas när det gäller parlamentets rättigheter .
Ändringsförslag 10 kan kommissionen , tyvärr , inte godta när det gäller tremånadersperioden och den mottagande medlemsstatens roll .
Kommissionen stöder i det avseendet ändringsförslag 22 , vilket jag redan påpekat .
Övriga ändringsförslag kan inte godtas .
Personligen känner jag sympati för namnet " EU-kort för tillhandahållande av tjänster " som föreslås i ändringsförslag 1 men Amsterdamfördraget tillåter inte det .
I ändringsförslag 18 hänvisas till direktiv 96 / 71 angående minimilöner som redan tillämpas , så det behövs ingen ändring .
Om kommissionen skulle godta ändringsförslag 17 så skulle det innebära att en enkel anmälningsplikt skulle gälla om inget giltigt kort lämnats .
Det är väl ändå i strid med intressena i samband med den allmänna ordningen i medlemsstaterna .
Ändringsförslag 19 är också oacceptabelt med hänsyn till mina beaktanden kring ändringsförslag 10 .
Kommissionen har samma ståndpunkt när det gäller liknande ändringsförslag till det andra förslaget .
Jag vill tillfoga att ändringsförslag 10 är helt godtagbart när det gäller det förslaget .
Med avseende på ändringsförslag 15 om definitionen av begreppet " egenföretagare " skall kommissionen , som jag redan sagt , se till att ta fram en nöjaktig lösning för att tillmötesgå de invändningar som rests .
Då övergår jag till Lord Inglewoods anmärkning .
Han hänvisade till de gränskontroller som finns med avseende på Förenade kungariket och jag skulle vilja säga att ingen medlemsstat , och alltså inte heller Förenade kungariket , har skyldighet att avskaffa kontrollerna vid de gränser som fortfarande finns .
Det gäller , som sagt , även för Belgien där den aspekten nyligen var aktuell .
Angående Karas anmärkning skulle jag vilja säga att jag fick intrycket att han talade om möjligheten att arbetstagare från Polen utnyttjas i hans land .
Kommissionen skulle vilja föreslå en lösning på det problemet varvid den lösningen skulle gälla för alla företag i Europeiska unionen som anställer personal från länder utanför EU .
Frågan är sedan om de två fallen skall behandlas lika .
Det är en fråga som jag tycker hör hemma i debatten om Europeiska unionens utvidgning och kanske inte i den här debatten .
För kommissionens räkning ställer jag mig gärna till Karas förfogande om han skulle vilja ha ytterligare information i denna mycket viktiga fråga .
Jag står alltså till förfogande .
Avslutningsvis skulle jag vilja tacka parlamentet för den mycket konstruktiva debatten om de viktigaste aspekterna av de här förslagen och speciellt naturligtvis den viktigaste föredraganden , Berger .
Tack så mycket , kommissionär Bolkestein .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.00 .
 
Förstainstansrätten Nästa punkt på föredragningslistan är betänkande ( A50003 / 2000 ) av Marinho för utskottet för rättsliga frågor och inre marknaden om I. förslaget till rådets beslut om ändring av beslut 88 / 591 / EKSG , EEG , Euratom om upprättandet av Europeiska gemenskapernas förstainstansrätt ( 5713 / 1999 - C5-0020 / 1999 - 1999 / 0803 ( CNS ) ) och II. förslaget till rådets beslut om ändring av beslut 88 / 591 / EKSG , EEG , Euratom om upprättandet av Europeiska gemenskapernas förstainstansrätt ( 9614 / 1999 - C5-0167 / 1999 - 1999 / 0805 ( CNS ) ) .
Herr talman !
Det är inte säkert att den framtida revideringen av fördragen under regeringskonferensen kommer att öppna dörrarna till en revidering av gemenskapens rättsordning .
Idén att ta med den här frågan i den dagordning som vi i dag diskuterar har stått fast sedan toppmötet i Helsingfors , den försvaras fortfarande av en del medlemsländer och hålls levande i Europaparlamentet , där utskottet för rättsliga frågor enligt min mening håller på att förbereda ett högkvalitativt uttalande om rättsreformens beskaffenhet och räckvidd .
Nästa gång parlamentet lägger fram ett betänkande om regeringskonferensens förberedelse så är jag övertygad om att man på grund av tre , som jag ser det , förenliga skäl med eftertryck kommer att ta upp frågan på nytt : Därför att rättvisa behöver skipas på kortare tid , därför att den rättsliga grunden för området för frihet , rättvisa och säkerhet måste skapas och till sist därför att sättet att se handel och ekonomi inom det europeiska området måste förändras genom att medborgarna övertygas om att de är en del av gemenskapsrätten som , baserad på en demokratisk lag och på domstolarna , respekterar de grundläggande etiska och juridiska värdena samt värnar om deras intressen , även om den nationella lagen inte är tillräcklig för att kunna garantera obegränsat medborgarskap .
Sanningen är att de förutsättningar som rättfärdigar en djupgående reform av gemenskapens rättssystem i dess helhet är också de som kan rättfärdiga en eventuell reform av Förstainstansrätten som vi i dag har uppe till behandling , men med en annan rättslig grund , det vill säga Amsterdamfördragets grund .
Det är i första hand två eller tre anledningar som legitimerar detta och som jag tänkte nämna : en bristande jämvikt mellan ett ökat antal rättsprocesser och den tekniska och mänskliga kapaciteten vid Luxemburgs domstolar , en rigorös skyldighet att erbjuda processuell flerspråkighet , ett korollarium till respekten för språk och nationella rättsliga traditioner , och till sist det faktum att domstolen - Förstainstansrätten - är enda instans för ekonomiska tvister där medborgare och företag kan anföra besvär mot myndighetsbeslut som påverkar dem .
Förslaget om att utöka antalet domare till 21 är därför helt och hållet berättigat , vilket till syvende och sist har att göra med domstolens effektivitet , samtidigt som man underlättar inrättandet av två extra salar för överläggning av information med vardera tre domare .
Den andra reformen har att göra med Förstainstansrättens utvidgade befogenheter , dit man hittills bara har kunnat kanalisera privatpersoners överklaganden och som nu också öppnas för medlemsstaternas besvärsskrifter .
Det som står på spel är ländernas möjlighet att överklaga ärenden som berör transportpolitik , konkurrensregler tillämpliga på företag , statligt stöd , åtgärder för handelsskydd , nyttjande av medel och andra åtgärdsprogram där hänsyn tas till beviljandet av finansiellt gemenskapsstöd , i första hand medel som berör unionens budgetmissbruk .
När möjligheten att överklaga till Förstainstansrätten öppnas för medlemsstaterna , där man nu kan processa om samma sak som en privatperson , kommer domstolen att få veta vilka överklaganden varje medlemsstat har gjort , vilket innebär att länderna och privatpersonerna blir jämlika i domstolens ögon .
Herr talman , man kan säga , menar några , att reformen är ytlig , men reformen är möjlig och grundar sig på normer som är tillämpliga i enlighet med Amsterdamfördraget .
I grund och botten är det ju faktiskt den som förutsågs och begärdes av gemenskapernas domstol , oberoende av regeringskonferensen och på grundval av nu gällande fördrag .
Eftersom kommissionens bifall var stort så lutar jag åt att parlamentet kommer att samtycka till de här två reformförslagen , ge domstolen sin röst och det enda som sedan fattas är att hoppas att också rådet gör detsamma .
Det är min slutgiltiga röst , måtte domstolen använda sin nya makt på bästa sätt , de nya befogenheter som parlamentet till sist gav den .
Herr talman !
Jag vill börja med att gratulera föredraganden till ett betänkande , som vid en första genomläsning endast ger intryck av att bekräfta och acceptera .
Bakom det här betänkandet döljer sig emellertid ett omfattande och effektivt arbete som redan har lett till vissa resultat : handlingens införlivande i det finska ordförandeskapets löfte den 7 december 1999 om att utvidga dagordningen för regeringskonferensen till att omfatta en undersökning av de framtida förändringarna av gemenskapens domstolars organisation , sammansättning och behörighet .
Därför vill jag framföra mitt erkännande av vice ordförande Marinhos insats .
Herr talman , en reform av gemenskapens rättsväsende har blivit en nödvändighet om man i framtiden skall kunna skipa rättvisa inom rimliga tidsramar , om Europeiska unionen i framtiden vill ha en rättskipning på samma nivå som det politiska projekt som vi har påbörjat .
I dag - och det säger jag med stolthet och glädje - har vi här i parlamentet haft ett ypperligt tillfälle att visa i vilken utsträckning vi européer anser att det politiska projektet är betydligt mer än den inre marknaden , ett projekt som i större utsträckning baserar sig på principer än på ekonomiska intressen .
För bakom principerna , herr talman , döljer sig alltid rättvisan .
Men justice delayed is justice denied ( att skjuta upp rättvisan är det samma som att neka den ) , och det är något vi bör fundera över .
Oroväckande uppgifter framkommer av det arbetsdokument som domstolen själv har förberett .
Mot bakgrund av detta är reformprojektet under föredragande av vice ordförande Marinho välkommet .
Denna lösning är ett lappverk , men även ett lappverk får duga , för vi kan för närvarande inte - något som han har påpekat - förvänta oss en stor reform av systemet på regeringskonferensen .
Vi måste komma med lösningar som , även om de är provisoriska , bidrar till en snabbare och effektivare rättskipning .
Det är två saker jag vill ta upp i det här inlägget , och som faller utanför själva betänkandet , på grund av den skyldighet som parlamentet enligt fördraget har att utarbeta ett kort och koncist betänkande utan någon fördjupning .
Det är två förslag från vice ordförande Marinho som , det vågar jag nog påstå , stöds av hela utskottet för rättsliga frågor och den inre marknaden .
Det första innebär att domarna i förstainstansrätten skall förses med ytterligare en référendaire .
Det andra är att översättningstjänsten vid förstainstansrätten skall skiljas från den vid domstolen .
I dagsläget måste förstainstansrätten vänta mycket länge på att få sina domar översatta .
Vi utgör en gemenskap , vars grundläggande princip enligt fördraget är en kulturell och språklig mångfald , och vi får under inga omständigheter överväga att avskaffa en sådan viktig möjlighet som att få ta del av en dom på det egna språket .
När vi ändå talar om regeringskonferensen , låt oss då tänka på två saker .
Det första gäller detta parlament .
Jag tror inte det skadar att vi insisterar på en större medverkan vad domstolen beträffar , och då även i utnämnandet av domarna .
Vi vill framför allt och i första hand att domstolens behörighet skall utvidgas samtidigt som förmågan att uppfylla sina skyldigheter , det vill säga dess resurser .
Vi vill att behörigheten skall utvidgas , i synnerhet vad gäller avdelning IV i EG-fördraget och avdelning VI i EU-fördraget , och att man i förbifarten undersöker vissa alternativ på dessa områden som är så utomordentligt viktiga för våra medborgare .
Då syftar jag åter igen på de uttalanden som vi har fått ta del av de senaste dagarna .
Herr talman !
Jag vill gratulera föredraganden och välkomna innehållet i detta betänkande .
Det har fått mig att tänka på två problem som jag har fått nyligen i mitt eget valdistrikt .
Båda gäller nära förestående avgörande i EG-domstolen .
Det första fallet gäller en stor hängbro och om brotullarna för den skall vara momspliktiga eller inte .
Beslutet skulle få enorma följder för vår lokala ekonomi .
Det andra fallet gäller en dam som skall pensioneras inom tretton veckor och som förtvivlat väntar på ett domstolsavgörande som allvarligt kommer att påverka hennes ekonomiska villkor som pensionär .
Detta är bara två exempel på verkliga vardagliga problem som förseningar i Europas rättssystem skapar .
Dessa förseningar kan innebära personliga svårigheter och även tragedier .
Med detta säger jag inte att alla våra egna nationella rättssystem fungerar perfekt men alltför ofta kan det hända att de väntar på ett förhandsavgörande från EG-domstolen .
Statistiken visar en oroande stigande trend i fråga om den tid som krävs för att hantera förhandsavgöranden .
Detta skall inte ses som kritik av domstolen eller dess personal utan snarare domstolens struktur och dess brist på resurser i en växande europeisk union .
Förslagen i detta betänkande är mycket välkomna som ett tillfälligt avhjälpande åtgärd , men Europa är en rättslig konstruktion och dess domstolar är avgörande för att allt skall fungera på vederbörligt sätt .
I avvaktan på den kommande utvidgningen måste regeringskonferensen ta itu med grundläggande reformer och omstrukturering av domstolssystemet .
I annat fall kommer vi alla , som valda representanter , att få ta emot mer och mer högljudda krav från våra medborgare då de inte får tillgång till snabba och effektiva rättssystem .
Herr talman , mina damer och herrar , kolleger !
Jag vill också tacka föredraganden för detta utmärkta betänkande .
Jag är också helt införstådd med hans slutsatser , där han särskilt föreslår att antalet rättssekreterare för domarna vid förstainstansrätten skall ökas och att förstainstansrätten skall ges en egen översättningstjänst .
Jag anser att detta faktiskt är nödvändigt , eftersom vi vid utskottets för rättsliga frågor besök i Luxemburg fick höra att , EG-domstolen , naturligtvis med naturnödvändighet , så att säga ofrånkomligt , har företräde framför förstainstansrätten vid utnyttjandet av den gemensamma översättningstjänsten , och att därför viktiga saker ofta inte kan behandlas tillräckligt vid förstainstansrätten .
Men jag anser också att reformerna måste gå längre än vad vi nu kommer att besluta om .
Jag tror att det exempelvis är värt att överväga att man på de områden , där redan domarkollegier , som liknar domstolar , i förväg fäller ett avgörande - jag vill bara nämna Alicante eller hur nu detta har planerats för den europeiska ämbetsmannalagen - i förekommande fall gör förstainstansrätten till sista instans , och här upprättar en avslutande behörighet .
Jag inser också att vi förmodligen måste göra något i samband med kommissionens tendenser att åternationalisera konkurrensavgöranden och lägga tillbaka dem på den nationella nivån .
Här förefaller det nödvändigt att överväga detta , eftersom dessa fall ju då inte längre skulle hamna hos förstainstansrätten , utan som förlagor till beslut vid EG-domstolen .
Vi bör överväga hur vi skall hantera denna situation .
Eventuellt bör det också finnas möjlighet att lämna förlagor till beslut i konkurrensärenden till den specialiserade avdelningen vid förstainstansrätten .
Dessutom måste man också överväga , om det är rätt - och vi har just haft fall , där ledamöter eller grupper har överklagat mot Europaparlamentet - att förstainstansrätten är ansvarig för sådana frågor , även om det egentligen handlar om författningsfrågor och dessa saker helt logiskt egentligt hör hemma hos EG-domstolen och mindre hos förstainstansrätten .
En sista punkt : Jag tror också att det behövs en demokratisk kontroll av OLAF .
För ögonblicket befinner sig OLAF i ett vakuum och kan göra vad den vill .
Jag anser att det är nödvändigt att OLAF kontrolleras av en domstol .
Den enda domstol som kan göra det på ett förnuftigt sätt skulle vara förstainstansrätten .
Också detta skulle vara en impuls för den fortsatta reformprocessen .
Herr talman !
Jag skulle vilja börja med att instämma med dem som gratulerade föredraganden för detta dokument .
Europeiska unionen är ett system grundat på lagar .
Den måste därför ha ett domstolsväsen för att genomdriva dessa lagar .
Om domstolarna dessutom inte kan klara av den arbetsmängd som läggs på dem på ett riktigt och snabbt sätt händer det som Palacio Vallelersundi redan påpekat , nämligen att försenad rättskipning blir samma som nekad rättskipning .
Domstolens bevis är att det händer nu och det pekar mot åtgärder som kan vidtas nu för att lindra problemet .
Men som Marinho påpekade , mer krävs , men det får vänta till regeringskonferensen .
I mitt eget land talas det mytiskt om de myllrande horderna av anonyma Brysselbyråkrater men man talar aldrig om antalet europeiska domare .
Det finns mindre än tre dussin i toppen på det europeiska rättskipningssystemet - knappast en överbemanning med tanke på deras ansvarsfulla uppgifter i hjärtat av det europeiska rättssystemet .
Hur stor deras betydelse är kan man se i de politiska följderna av förseningen med att lösa den mycket viktiga engelsk-franska tvisten om brittiskt nötkött som har skapat så mycket ilska i mitt land och sådan besvikelse över unionens handläggning av domstolstvister .
Detta har förvärrats , något som några av mina rådgivare anser , av procedurreglerna i de franska domstolarna som gör det nästan omöjligt för icke franska medborgare att öppna process mot den franska regeringen .
Det uppfattas faktiskt som omöjligt .
Detta kontrasterar mycket ofördelaktigt mot Förenade kungarikets domstolar där spanska fiskare framgångsrikt lyckades väcka åtal mot Förenade kungarikets regering under mycket jämförbara förhållanden .
Vad som händer i Frankrike , herr talman , verkar vid första anblicken vara ett fall av diskriminering mot övriga EU-medborgare på grund av nationalitet och därmed bryta mot fördragen .
Jag skulle därför vilja be kommissionären , som var vänlig nog att kommentera mina inlägg i den tidigare debatten , att undersöka detta och meddela resultaten till parlamentet och mig .
Jag skulle vara tacksam om kommissionären i sin slutkommentar kan bekräfta att han kommer att göra detta . .
( NL ) Herr talman !
Å kommissionsordförande Prodis vägnar skulle jag gärna vilja svara så här .
Kommissionen noterar den ståndpunkt som Europaparlamentet i dag intagit angående domstolens och förstainstansrättens begäran om att å ena sidan till förstainstansrätten överlåta den bedömning av vissa överklaganden som domstolen nu har ensam behörighet för och å andra sidan öka antalet ledamöter i förstainstansrätten .
Jag skulle vilja tillfoga att jag för kommissionens räkning med stort intresse lyssnat till de anföranden som hållits här alldeles nyss och att jag mycket väl begriper den oro som ligger till grund för dessa anföranden .
Den oron är berättigad .
Det har flera gånger sagts att justice delayed is justice denied .
Kommissionen begriper den inställningen .
Mot bakgrund av den insikten skulle jag vilja fortsätta mitt svar på följande sätt .
Som parlamentet vet så är kommissionen övertygad om att gemenskapens rättsinstanser utan en grundlig reform löper risken att på kort sikt inte längre kunna utföra sina uppdrag inom rimliga tidsfrister .
Kommissionen har därför också rådfrågat en expertgrupp om de reformer som skulle kunna genomföras för att domstolen och förstainstansrätten skall behålla kvaliteten och koherensen i sina domslut under kommande decennier .
Kommissionen känner till förstainstansrättens begäran om personalförstärkning men för ögonblicket anser kommissionen att den föreslagna överföringen av behörigheter skall betraktas i ljuset av den undersökning som jag nyss nämnde och kommissionen skall lämna sitt yttrande om domstolens och förstainstansrättens begäran i ljuset av den undersökningen , alltså så snabbt som möjligt efter att undersökningen slutförts .
Tack , herr kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11 .
 
Exceptionellt finansiellt stöd till Kosovo Nästa punkt på föredragningslistan är betänkande ( A5-0022 / 2000 ) av Brok för utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik om rådets förslag till beslut om exceptionellt finansiellt stöd till Kosovo ( KOM ( 1999 ) 0598 - C5-0045 / 00 - 1999 / 0240 ( CNS ) ) .
Jag har fått veta att vår föredragande är försenad några minuter .
Jag föreslår att vi inleder debatten omedelbart .
Föredraganden är på väg hit och kommer att tala så fort han anlänt .
Jag lämnar därför ordet till Bourlanges i hans egenskap av föredragande av yttrandet från budgetutskottet .
Herr talman !
Denna fråga är viktig och brådskande och parlamentet , som ombetts av kommissionen att snabbt uttala sig , gör det också , för man skall veta att i dag dör män och kvinnor i Kosovo , helt enkelt för att det är 25 grader kallt , att dessa människor utför ett enormt arbete för att garantera ett minimum av underhåll och att de inte får betalt .
Vi har därför mottagit en begäran om brådskande förfarande som vi beviljar .
Man ber oss om 35 miljoner euro .
Vi är överens om att ge ut dem och vi ber kommissionen att visa prov på stor vaksamhet så att beloppen verkligen betalas ut så fort som möjligt när beslutet väl har fattats .
Det är fråga om makroekonomiskt stöd .
Det orsakar reaktioner på vissa ställen eftersom de liberala idealen inte respekteras som består i att ingripa ekonomiskt för att stödja en administration .
Det är inte vår uppfattning .
Vår uppfattning är att det är grundläggande att bidra till att inrätta en administration i Kosovo och att det inte alls är absurt att direkt bidra till att betala de offentliga tjänstemännen i denna region .
Det skulle för övrigt ha varit något mycket användbart som vi skulle ha kunnat göra i Ryssland under hela 90-talet för att undvika denna stats upplösning .
Det andra stora problemet är att man vänt sig till oss , givarna har gjort åtaganden men vi är uppenbarligen de enda som betalar .
De andra betalar inte .
Vi kräver att denna unilaterala situation skall upphöra när det gäller att begära ekonomisk hjälp .
Vi önskar att kommissionen gör utfästelser när det gäller våra ändringsförslag i det hänseendet .
Vi vill knyta beviljandet av hela stödet till mobiliseringen av pengar som övriga givare är skyldiga .
Inte för att begränsa , för att knussla med vårt ekonomiska stöd till Kosovo utan tvärtom för att se till att vårt stöd kommer utöver det från övriga givare .
Ur den synvinkeln är den bestämmelse som föreslås en bestämmelse om stöd i två etapper och den andra bör frigöras när givarna visat att de är intresserade .
Avslutningsvis ställer vi tre frågor till kommissionen i detta hänseende : för det första måste den på ett regelbundet sätt ge oss förteckningen och beloppen när det gäller bidrag från övriga givare .
Vi vill veta vad de övriga betalar när vi betalar .
För det andra vill vi ha en exakt lägesrapport över anbudsinfordran och deras åtagandetakt .
Man sade oss under budgetförfarandet att det var brådskande att rösta för pengarna till Kosovo och enligt den information vi förfogar över har hittills ingen anbudsinfordran offentliggjorts eller inletts .
Det är allvarligt eftersom det försenar hela återuppbyggnaden av Kosovo .
Avslutningsvis , och det är konsekvensen av vad jag just sagt , vill vi att kommissionen mycket regelbundet , varje månad , informerar budgetutskottet om läget för verkställandet av utgifterna .
Vi har papper från kommissionen där man talar om bestämda åtaganden .
Vi behöver inga bestämda åtaganden , vi behöver åtaganden helt enkelt och vi behöver veta vad som verkligen betalats och framför allt vad som inte betalats .
Kosovo har lidit alltför mycket av försenade betalningar .
Herr talman !
När vi i dag talar om Kosovo , vilket vi ju ofta har gjort , bör vi också någon gång avlägga räkenskap om vad som redan har gjorts i Kosovo , eller om det över huvud taget redan gjorts något .
Jag anser att man redan har tagit några små steg på vägen mot en normalitet , och man skulle åtminstone vilja räkna upp dem inom ramen för en sådan debatt .
Det finns från och med den 9 februari ett s.k. interimsråd - man kallar det Kosovo Transitional Council - , där både de politiska partierna , minoriteterna och the civil society är representerade , och som skall fungera ungefär som ett interimsparlament .
Det är bra , det välkomnar vi , men jag tror att man också måste ge dem ett instrument i handen och en strategiplanering för det som de egentligen bör förbereda , ty i höst planerar man att hålla val .
Ingen vet riktigt vad dessa val skall leda till , och vilket parlament som skall bildas .
Ingen vet vilka befogenheter detta parlament sedan skall ha gentemot UNMIK .
Det betyder att det finns många svårbedömbara saker som vi inte informeras om och som andra förmodligen inte heller kan riktigt förstå .
Just albanerna , som nu integreras i detta interimsråd , borde egentligen få en något bättre uppfattning om vad som väntar dem .
Vid sidan av det ekonomiska arbetet , vid sidan av återuppbyggnaden , måste man ovillkorligen också tänka på hur man skall åstadkomma någon samexistens mellan serber , albaner och andra minoriteter - exempelvis också zigenarna - så att det , på vägen till samexistens , någon gång i en nära framtid förhoppningsvis kan äga rum en försoning .
Jag vill än en gång räkna upp vad det redan finns av faktiska saker som vi kan glädja oss åt .
När det gäller förvaltningen finns det nu 34 skatteinspektörer .
Det är bra !
Människorna uppmanas nu också att betala sina skatter även där , ty på sikt kan det ju inte gå an att alla bara är beroende av EU : s och andra givares portmonnäer ; en del måste man även på detta område åstadkomma på egen hand .
Det kan dessutom fastslås att av 19 departement har redan 4 en administrativ ledning , vilket också är ett framsteg jämfört med vad vi tidigare haft där .
Vi har dessutom något som är mycket viktigt för den rättsstat som vi ju vill bygga upp .
Vi har 130 domare och åklagare , som nu har avlagt eden , och som kan ta upp sitt arbete för att skipa rätt , för att också litet grand berika toleranskulturen där en aning och naturligtvis också åtminstone komma förbrytelserna på spåren och då också kunna döma .
Det som också är bra , det vill jag erinra om , är det faktum att den gamla UCK nu är integrerad i återuppbyggnaden av detta land .
Jag tror att det är bra .
Jag ansluter mig helt och fullt till det som budgetutskottet har sagt i fråga om finansieringen , och jag anser att vi måste erinra kommissionen om att den verkligen måste insistera på att andra givare äntligen betalar sin andel .
EU-kommissionen kan inte betala för allting .
Den är där nere ansvarig för återuppbyggnaden , den är ansvarig för den fjärde pelaren , men den kan inte också alltid betala Kouchners löpande kostnader .
Det kan man göra en eller ett par gånger , men jag tror att FN : s givare också måste bidra till det , och där finns det ett mycket stort hål , som inte är fyllt , och som vi inte kan fylla .
Vi har en stor uppgift i återuppbyggnaden , det är vår uppgift , och vi bedöms efter hur vi utför denna uppgift !
Herr talman !
Jag vill göra några preciseringar .
Risken i en debatt är alltid att vi som medverkar upprepar oss för mycket .
Men jag skall koncentrera mig på fyra punkter .
Till att börja med vill jag fastslå att unionen är den största bidragsgivaren till återuppbyggnaden av Kosovo .
Och till Albright kan jag säga att detta har stått i tidningen på senare tid , och siffrorna ljuger inte .
Detta råder det ingen tvekan om , även om man kunde önska att det inte vore fallet .
Unionen har beslutat att bidra med ytterligare 35 miljoner euro i makrofinansiellt stöd till återuppbyggandet av Kosovo , mot bakgrund av en rapport från FMI där man uppskattar att återuppbyggandet kräver ytterligare 115 miljoner .
Jag vill nämna för Pack att jag med henne är helt överens om att kommissionen måste uppmana de övriga bidragsgivarna att uppfylla sina löften .
Dessutom vill jag ge uttryck för min oro - en mycket stark sådan - över vissa ministrars uttalanden på det senaste Ekofin-rådet , som visar att man vill att en av det portugisiska ordförandeskapets prioriteringar skall vara att den budgetplan som man enades om i Berlin under inga omständigheter ändras .
Detta innebär ett ifrågasättande av det avtal som parlamentet med stora svårigheter lyckades uppnå med rådet i december , enligt vilket man , när kommissionen lägger fram ett flerårigt program för återuppbyggandet , skall vidta en granskning av budgetplanen .
Därför vill jag uppmana dessa ministrar att inte ifrågasätta det avtal som var så svårt att uppnå .
Jag vill be kommissionen , och det gläder mig att kommissionär Solbes är här i kväll , att i god tid lägga fram detta fleråriga finansieringsprogram , med tillhörande rapport , enligt parlamentets begäran , så att det kan beaktas i framtagandet av budgetförslaget till nästa budget , i överensstämmelse med det som vi har blivit lovade .
Slutligen vill jag poängtera att vi även om vi nu har kommit överens om 35 miljoner , vet att det bara är en droppe i havet och att det inte är tillräckligt , och därför måste vi så snart som möjligt uppnå en överenskommelse om ett flerårigt program för det så nödvändiga återuppbyggandet av Kosovo .
Herr talman , kolleger !
Jag ber er ursäkta att jag är försenad , men i dag är tyvärr denna andra politiska fråga fortfarande på föredragningslistan .
Utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik rekommenderar att ni lösgör dessa 35 miljoner euro , och den rekommendationen ger man eftersom dessa pengar verkligen kan komma de drabbade människorna till godo .
Det vi är kritiska till är inte så graverande att vi inte vill hjälpa människorna där nere .
Men det betyder inte att vi glömmer bort kritiken .
Vi skulle naturligtvis redan ha kommit mycket längre i vårt förfarande om rådets förvaltning inte hade glömt bort att på ett tidigt stadium informera Europaparlamentet och officiellt lämna information till det .
Endast på så sätt hade vi kunnat genomföra ett verkligt förnuftigt , djupgående samråd i saken .
Jag ber förvaltningen att se till att detta inte kan hända i framtiden .
Endast för de drabbade människornas skull är vi beredda att bortse från det och dra konsekvenserna av det .
Men vi måste se till att vi här inför bestämda villkor .
Ett villkor är att pengarna ges dit där de kommer att användas på ett klokt sätt , och inte till dem som möjligen kan använda pengarna för att tjäna andra syften , dvs. dessa pengar bör verkligen gå in i Kouchners ansvarsområde och inte till andra områden .
För det andra : Även om kommissionen och rådet här intar en annan ståndpunkt , eftersom de där ser realistiska problem , anser vi att de andra givarna också måste uppfylla de åtaganden som de har ingått .
Detta är en mission som står under FN : s ansvarsområde , och det får inte vara så att enbart Europeiska unionen uppfyller sina förpliktelser !
De andra givarländerna måste uppfylla sina förpliktelser på samma sätt under denna tidsrymd till gagn för de drabbade människorna .
Detta får mig att anse att vi i framtiden rent allmänt måste befatta oss mycket intensivare med denna fråga , och inte bara när det gäller detta konkreta projekt , utan hela utvecklingen i Sydosteuropa , och den hjälp som lämnas där .
Detta är återigen ett exempel för att Europeiska unionen är beredd att hjälpa till att ge pengar , men att den politiska ledningen inte är enhetlig .
Vi har så många samordnare , som är ansvariga inför så många arbetsgivare , att vi snart måste tillsätta en samordnare för samordnarna .
Men det kanske vore bättre om de ansvariga instanserna i Europeiska unionen och de andra institutionerna , från OSSE till Förenta nationerna - skulle sätta sig ned för att införa ett enhetligt , samordnat förfarande , och granska hur man verkligen kan hjälpa människorna där .
Jag vet att man inom kommissionen intensivt funderar över hur man skall uppnå detta , men om Europeiska unionen bidrar med den största delen , då skall den också ha hand om ledningen där och sedan sköta det på ett enhetligt sätt , så att människorna verkligen blir hjälpta .
Det är ingen mening med att vi här snarast har en konkurrens mellan de olika internationella inrättningarna och sammanslutningarna , i stället för att kraften verkligen utnyttjas för att hjälpa människorna på platsen !
När jag ser att givarkonferensen för stabilitetspakten hela tiden skjuts upp , nu till slutet av mars , och att ingen vet vilka projekt som verkligen ligger bakom , när man inte kan överblicka på vilket vis det verkligen kan genomföras , och det hela tiden ges nya presskonferenser , då verkar detta inte vara rätt sätt att skapa fred och försoning mellan människorna i denna del av Europa !
Av den anledningen , kära kommission , kära ordförandeskap i rådet , vill vi också ta detta till anledning för att uppmana er att gripa detta politiska initiativ , så att vi inte åter hamnar i en sådan nödsituation att vi i slutet av en månad måste ordna upp betalningsförmågan , utan att det därmed kan ställas upp en långfristig strategi för hjälpen i denna region , och jag hoppas att ni då äntligen kan uppfylla era politiska förpliktelser , och att det inte fortsätter så som vi har upplevt det under de senaste månaderna !
Herr talman !
När alliansen engagerade sig i Kosovo var det med målsättningen att i denna provins återupprätta villkor som gör det möjligt för dem som så vill att stanna kvar , återvända till sina rötter och till sin egen kultur .
Om alliansen i dag är närvarande på fältet är det med samma målsättning .
I förrgår lyssnade jag med tillfredsställelse till en intervju med en befälhavare i Kfor som berättade att saker och ting började fungera bättre i Kosovo och att normerna för brottsligheten återgått till en acceptabel nivå , framför allt när det gäller säkerhet .
De som befinner sig på fältet för att företräda Europa och fortsätta med dessa målsättningar , och jag tänker särskilt på den särskilda representanten för Förenta nationernas generalsekreterare , är nära att ge upp , just på grund av det faktum att situationen förbättrats och man talar mindre om Kosovo , och att det därför är mindre uppenbart hur brådskande hjälpen är som behöver beviljas .
Vi måste arbeta för att se till att epoken med kommers ersätter den med krigsherrarna , i denna provins liksom i hela Balkan i allmänhet .
Det ekonomiska stödet är i det hänseendet en beståndsdel som förvisso är grundläggande när det gäller möjligheter till åtgärder för dem som befinner sig på fältet .
Jag upprepar här Doris Packs uttalande och jag betonar att vi i Europaparlamentet måste ta vårt ansvar i detta hänseende , men vi skall naturligtvis se till att vi inte är ensamma om det .
Herr talman , herr kommissionär , mina damer och herrar !
Först vill jag tacka föredraganden , kollegan Brok , så hjärtligt för hans betänkande .
Om rådet hade arbetat så snabbt som kollegan Brok gjort , då skulle vi i själva verket ha kommit mycket längre .
Rådets försummelse kan man här verkligen beklaga !
Föredraganden och betänkandet utgår helt riktigt från att vi bör och måste lämna snabb hjälp , men de utgår också helt riktigt från att vi inte skall lämna obegränsad eller godtycklig hjälp .
Här vill jag i synnerhet hänvisa till ändringsförslag 5 , där det helt klart fastslås att man med hjälp av medlen från det särskilda ekonomiska stödet uteslutande kan och får finansiera sådana budgetbehov i Kosovo , som uppstår i offentliga / halvoffentliga , kommunala och övriga förvaltningar och institutioner , som direkt eller indirekt kontrolleras av UNMIK .
Det måste stå klart , herr kommissionär , att vi stöder UNMIK , vi stöder de institutioner som inrättats av Förenta nationerna , i synnerhet naturligtvis pelare 4 , och det går inte an att vi stöder parallella strukturer som har bildats i Kosovo och fortfarande finns kvar där .
Vad skall nu göras med dessa pengar ?
Jag vill särskilt hänvisa till de mänskliga rättigheterna .
Västmakterna har i Kosovo kämpat för de mänskliga rättigheterna .
Vad sker i dag i Kosovo ?
Den stora aktionen för att driva bort serberna kunde stoppas , men nästan dagligen sker det oacceptabla saker , människor dödas , människor hindras att leva där , och att leva på sitt vis .
Dagligen sker det angrepp på serber , på zigenare , på bosnier , men det sker också fortfarande angrepp på albaner .
Jag blev förskräckt när jag läste betänkandet , om det nu stämmer att en albansk läkare , som säkerligen med stora svårigheter arbetat i sjukhuset i Mitrovic i den serbiska delen , slutligen gav upp att arbeta för sin befolkning i detta sjukhus , eftersom han hela tiden hotades till livet .
Detta är händelser och situationer som vi inte kan acceptera .
Jag har hört - om det stämmer vet jag inte - att serberna fortfarande rent av driver en gruva i Kosovo , i den serbiska delen .
Det finns åtminstone rykten om att serbisk milis fortfarande är aktiv .
För mig är det betydelselöst om det är en serb , en zigenare , en bosnier eller en alban som hotas eller dödas i Kosovo .
För mig är det betydelselöst vem som arbetar på att dela Kosovo .
Det som är avgörande för mig är att de organ som finansieras av oss uppnår det som vi vill uppnå , nämligen ett multietniskt Kosovo , ett liv sida vid sida i Kosovo .
Vi behöver mer polis , det finns absolut inte tillräckligt med polis .
Vi behöver ett oberoende rättsväsende - det är säkert svårt att bygga upp - och vi behöver också anslag för den höge kommissionären för de mänskliga rättigheterna .
Allt detta måste ske , och det måste ske snabbt .
Om vi inte snabbt lämnar hjälp , då kommer situationen att förvärras , och det kan uppstå nya konflikter och krissituationer .
Därför anser jag att det var rätt att vi handlade snabbt , att vi bekräftade att det var brådskande , och att vi ställer pengarna till förfogande .
Men vi vill se vad som görs , och vi vill också se resultat i Kosovo , och jag ber kommissionen att se till att dessa pengar också används med framgång , i synnerhet för att bygga ut polisväsendet och rättsväsendet . - Herr talman !
Till en början ett stort tack till ledamöterna , och i synnerhet till föredraganden , för den snabba behandlingen av denna fråga .
Det kommer utan tvivel göra det möjligt för oss att snabbt frigöra medel till Kosovo och ta oss an de orosmoment som både Swoboda och Pack har påtalat .
I den här kvällens debatt tycker jag mig märka tre starka orosmoment .
För det första är det sant att vi , även om det har skett stora framsteg , och där kan nämnas tullförvaltningen , bankförvaltningen och skatteförvaltningen , måste fortsätta framåt .
Framåt mot en finansiering av vad ?
Där har vi den första punkten där det råder en viss oenighet .
Ni föreslår i ett av era ändringsförslag att enheterna som är föremål för unionens finansieringsbidrag skall begränsas mer .
Till exempel i ändringsförslag 3 och 5 .
Emellertid bör man , enligt vår uppfattning , i båda avseendena lämna större handlingsutrymme åt Förenta nationernas förvaltning som känner till förhållandena på platsen bättre än vi .
Vi anser att det skulle innebära stora praktiska svårigheter att redan på förhand definiera vart resurserna skall gå .
Vi måste utan att tveka förlita oss på dem som där på plats , på ett bättre sätt än vi , kan fatta vissa beslut .
Det andra orosmoment som jag har förstått att vissa av er känner av - det lades till att börja med fram av Bourlanges , och det har upprepats av andra - gäller det som händer med övriga bidragsgivare .
Är det så att kommissionen gör en överdriven insats , medan de övriga struntar i att samarbeta ?
Vissa av ändringsförslagen i ert betänkande pekar i den riktningen .
Till exempel ändringsförslag 1,2 och 4 .
Jag kan tala om för Bourlanges och för dem som har lagt fram denna fråga , att det främsta problemet inte gäller tanken som sådan , som vi är helt eniga i .
Det främsta problemet är att fördelningen av bördan mellan de olika bidragsgivarna för närvarande har fastställts - och det är sant - i uttalandena av high level steering group , men det stämmer också att de saknar juridiskt värde , att det endast rör sig om ett politiskt åtagande .
Det är anledningen till att vi ber att ändringsförslag 1 , och vi har meddelat Brok detta , med bibehållen andemening skall formuleras på ett annat sätt så att det inte innehåller några villkor för tilldelningen av gemenskapens resurser .
Det samma gäller ändringsförslag 2 , som vi också finner godtagbart om det bara justeras något , eftersom vi anser att idén vad det finansiella stödet beträffar i sig är korrekt .
Ungefär samma sak gäller ändringsförslag 4 .
I denna konkreta fråga är det möjligt att vi har ett mer positivt besked till Bourlanges .
Rådet är redan vidtalat , så att det skall låta sitt beslut omfatta ett uttalande av kommissionen där detta villkor fastslås .
Det vi föreslår är närmare bestämt , vad det andra bidraget beträffar , att det exakta totalbeloppet och tidpunkten för den andra delutbetalningen skall avgöras med hänsyn till Kosovos externa finansiella behov och stödet från övriga bilaterala bidragsgivare .
Vi fastslår med andra ord inget villkor , eller vi tror att det är mer effektivt att inte fastslå något villkor från början , och ändå gör vi det beträffande detta eventuella frigörande av den andra delutbetalningen .
På det viset kommer vi inte att ha några problem med att agera omedelbart , vi skapar inga problem för befolkningen i Kosovo , men däremot tvingar vi de övriga bidragsgivarna att genomföra sina finansiella insatser på samma sätt som vi gör .
Ett tredje problem har påtalats av Dührkop beträffande de fleråriga programmen .
Jag kan påminna om att projekten är fleråriga .
I programmen måste man givetvis ta hänsyn till det årliga budgetstödet .
Till slut vill jag kommentera de önskemål som har framförts om ytterligare information .
Å ena sidan har man bett oss underlätta utvecklingen av anbudsförfarandet för parlamentet , och på den punkten kan jag tala om för er att kommissionen redan förra veckan hade tillfälle att ge parlamentets budgetutskott en lägesrapport om de kontrakt och betalningar som har utförts sedan task force började fungera i Kosovo .
Kommissionen kan lova att även framöver regelbundet informera parlamentet om de anbudsförfaranden som offentliggörs .
Vår önskan är att detta även läggs ut på Internet , så att största möjliga insyn ges i denna konkreta fråga .
En annan sak jag vill kommentera är övrig information som kan vara av betydelse för parlamentet vad gäller det makroekonomiska stödet .
I det avseendet kan jag även meddela att kommissionen är villig att regelbundet informera ordförandena i de olika parlamentsutskott som är involverade i frågan , under konfidentiella former om den information som ges förutsätter detta , samt utifrån de olika planer som tillämpas för de makroekonomiska stödåtgärderna .
Ett stort tack till alla ledamöter , och jag hoppas att vi i och med rådets slutgiltiga beslut kan få loss dessa medel och förverkliga ett positivt stöd som gör det möjligt för oss att fortsätta med de viktiga insatser som görs i Kosovo från olika håll för att uppnå den situation som vi alla önskar med en ökad förståelse och fred .
Herr talman !
Jag gläds åt att åsikterna från parlamentet , särskilt budgetutskottet , och kommissionen är så samstämmiga , och vi försäkrar att för vår del kommer vi alltid att troget hjälpa kommissionen att genomföra sin uppgift .
Jag känner ändå en viss oro när jag lyssnar till kommissionären jämfört med de åtaganden som gjorts av enheterna inom budgetutskottet .
Det beslutades tydligt - jag säger inte att det var bra eller dåligt , men det var ett avtal - det beslutades tydligt mellan kommissionens enheter och budgetutskottet att man var överens om ändringsförslag 4 och 7 , dvs. man var överens om idén att knyta mobiliseringen , genomförandet , av den andra delen av det makroekonomiska stödet till respekten för de åtaganden som tidigare gjorts av givarna .
Men jag tyckte mig förstå när jag lyssnade till Solbes att detta åtagande skulle ske på ett diskret sätt .
Herr kommissionär !
Ett avtal är ett avtal .
Ja eller nej , bekräftar ni det godkännande som gjorts av era enheter i budgetutskottet eller släpper ni detta villkorande , vilket skulle innebära att ni bryter ett åtagande mot oss ? .
( FR ) Nej , herr Bourlanges , jag tror att det handlar om ett sakproblem .
Problemet är : hur skall vi styra den kompromiss vi accepterat .
Vad jag föreslog er , vad jag säger igen , är att kommissionen skall göra ett uttalande , i rådets beslut , i följande riktning : Det exakta beloppet och tidpunkten för att inleda den andra delen kommer i sinom tid att beslutas med hänsyn till utvecklingen av Kosovos yttre ekonomiska behov och bidrag från andra bilaterala givare .
Därför anser vi att vi fullständigt respekterar det som vi kommit överens om .
Jag begär bara att kommissionen skall informera budgetutskottet innan den andra delen genomförs . .
( FR ) Jag instämmer helt , och det kommer vi att göra .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11 .
 
Altener Nästa punkt på föredragningslistan är betänkande ( A5-0011 / 2000 ) av Langen om förlikningskommitténs gemensamma utkast till parlamentets och rådets beslut om ett flerårigt program för främjande av förnybara energikällor inom gemenskapen - Altener ( C5-0333 / 1999 - 1997 / 0370 ( COD ) ) Herr talman !
Jag tackar Langen - även om han inte själv är närvarande här - för det arbete som han lagt ner för att driva igenom programmet såväl i parlamentet som i rådet .
Projektet har varit långvarigt och besvärligt .
Man måste även i fortsättningen satsa särskilt mycket på sådan forskning som kartlägger användningen av förnybara energikällor .
Även om det nya direktivet innehåller mycket gott är det dock också behäftat med brister .
Ett exempel på detta är torven .
Torv får inte placeras i samma grupp som fossila bränslen .
Kan man inte direkt klassificera torven som en förnybar , icke-fossil energikälla måste man särskilt med tanke på miljöbeskattningen definiera en egen klass för den .
Det är inte rättvist att torven värderas på samma sätt som exempelvis stenkolen .
Utvecklingen av förnybara energikällor är en dellösning för att avskaffa unionens beroende av importerad energi .
Forskningen är av speciellt stor betydelse också med tanke på EU : s nästa utvidgningsrunda .
Beroendet av importerad energi berör allra värst just flera östeuropeiska länder vars ekonomiska struktur fortfarande lider av det beroende av rysk energi som skapades under sovjettiden .
EU måste hålla fast vid Kyotos klimatprotokoll .
Vi är ju alla bekymrade över miljön och våra barns framtid .
De förnybara energikällornas andel av den totala energiproduktionen måste ökas , men det måste också göras med förnuft .
Vi måste komma ihåg att vi inte på länge än kan bygga vår grundläggande energiproduktion på förnybara energikällor .
Där behövs energi som skonar klimatet , kärnkraft . .
( DE ) Herr talman !
Jag ber om överseende med att jag kommer litet sent , eftersom det hela ändå har förlöpt något snabbare än förväntat .
Jag tackar kollegan för att hon hoppade in i mitt ställe .
Hon har ju redan sagt något om programmen Altener och Save .
Vi har här slutuppgörelsen för ett förlikningsförfarande om åtgärder inom energiområdet för perioden 1998 - 2002 .
Altener behandlar där det viktigaste området beträffande de förnybara energikällorna .
Därigenom skall det skapas nödvändiga förutsättningar för att genomföra en handlingsplan på detta område , och i synnerhet skall det ges stimulans till privata och offentliga investeringar i produktion och utnyttjande av förnybara energikällor .
Eftersom det löpande programmet löpte ut i slutet av förra året och rådet inte godtog de ändringar som parlamentet beslutat om , måste förlikningskommittén träda i funktion .
Det är ganska förvånande att se hur envist medlemsstaterna i rådet försökt värja sig mot detta program för alternativa energikällor och mot rimliga anslag för detta .
Men jag måste också säga att den finske rådsordföranden var mer eller mindre oförmögen att agera så länge som medlemsstaterna blockerade den nödvändiga höjningen av dessa anslag .
Det ursprungliga förslaget om 81,1 miljoner euro , som föreslagits av kommissionen , sänktes ensidigt och utan motivering av rådet till 74 miljoner euro .
Det var därför bara följdriktigt att parlamentet krävde att det ursprungliga förslaget till anslag åter skulle läggas in .
Vid sidan av hur programmet skulle finansieras tvistade parlamentet och rådet också om vissa andra punkter .
Inom ramen för förlikningsförfarandet kunde man på väsentliga punkter , som krävts av oss , uppnå enighet med rådet , till exempel också undersökningen av möjligheten att öppna Altener-programmet för de associerade Medelhavsländerna med anledning av nästa revidering av detta program .
Till detta kommer rådet - det har man försäkrat oss - att i Europeiska gemenskapernas officiella tidning offentliggöra ett uttalande .
Med tanke på den ekonomiska ramen skulle rådet , genom att tydligt reducera sitt ursprungliga förslag , nästan ha äventyrat möjligheten att fortsätta med programmet .
För parlamentets delegation till förlikningskommittén handlade det om att fortsätta med innehållet i ett klokt program .
Därför röstade vi till slut för kompromissen , även om vi inte var fullt tillfreds med den .
Vi accepterade att medlen höjs till 77 miljoner euro .
Det är ett acceptabelt , om än inte helt tillfredsställande resultat .
Vi beslöt oss för denna kompromiss för att inte äventyra möjligheten att fortsätta programmet .
Utan förstärkta ansträngningar från medlemsstaterna förefaller det dock inte möjligt att uppnå målet att år 2010 täcka 15 procent av det totala behovet av energiförsörjning när det gäller primärenergi med hjälp av förnybara energikällor .
På så sätt garanteras det att ett miljö- och ekonomipolitiskt viktigt EU-program fortsätter , som bidrar till att begränsa koldioxidutsläppen , öka andelen förnybara energikällor i energibalansen , minska beroendet av energiimport , säkra försörjningen och hålla samman den lokala och regionala utvecklingen .
Men det räcker naturligtvis inte , utan det måste också göras väldiga ansträngningar från medlemsstaternas sida .
Förlikningskommittén antog den 9 december förra året den slutgiltiga texten för programmet och jämnade därmed vägen för att man för alternativa energikällor även i framtiden skall främja undersökningar och åtgärder för att exploatera potentialen med förnybara energikällor .
Dessutom garanteras det , genom att Altener-programmet fortsätter , att man kan stödja och genomföra pilotåtgärder för att skapa och bygga ut infrastrukturer , förmedla kunskap och vidta riktade åtgärder för att underlätta för förnybara energikällor att bli genomförbara och göra sig gällande på marknaden .
Detta är särskilt möjligt när det gäller jordvärme , vindenergi , mindre vattenkraftverk , passivt och aktivt utnyttjande av solenergi i byggnader och användning av biomassa .
Vi kan på dessa områden se hur nödvändigt och viktigt det är att även i fortsättningen ställa en förnuftig ram för stödåtgärder till förfogande för alternativa energikällor inom Europa .
Jag vill i synnerhet tacka kommissionen och den ansvariga kommissionären , de Palacio , för att hon stött parlamentets ståndpunkt .
Europaparlamentet har lyckats finna en förnuftig kompromiss och ändra rådets gemensamma ståndpunkt .
Jag vore tacksam om kollegerna kunde godkänna förlikningskommitténs resultat .
Herr talman !
Å PSE-gruppens vägnar är jag positiv till att vi har kommit fram till ett resultat i förlikningsförfarandet beträffande Altener II-programmet .
Men först vill jag tacka föredraganden , kollegan Langen , för hans verkligt bra arbete med detta betänkande .
Jag vill också tacka ledaren för delegationen till förlikningskommittén , kollegan Provan .
Ty som Langen just sade var det verkligen en hård kamp i förlikningskommittén .
Men vi kan i dag se att resultatet av förlikningen också absolut mycket tydligt visar vad Europaparlamentet förmår .
Langen påpekade att en rad punkter beträffande innehållet och krav från parlamentet införlivats , och när det gällde den viktigaste konflikten med rådet , anslagen till detta fleråriga program för att främja de förnybara energikällorna i gemenskapen , kunde vi - det har redan sagts - enas med rådet någonstans på mitten .
Det är inte tillfredsställande , det vill jag också säga helt klart .
Men vi har gått med på denna kompromiss , eftersom det var viktigt för oss att detta program nu verkligen kan startas mycket snabbt .
Ty under de närmaste åren skall andelen förnybara energikällor fördubblas till minst 12 procents andel av energiförbrukningen .
Det är Europeiska unionens uttalade mål .
Där har Altener-programmet verkligen en nyckelroll , som enda EU-program med den uteslutande målsättningen att främja förnybara energikällor .
Med detta nya femårsprogram måste dels åtgärderna från Altener I-programmet utökas .
Hit hör bland annat fördjupningen av informations- och erfarenhetsutbytet mellan aktörerna på området med alternativa energikällor , bland annat utbyggnad av lokala och regionala energiagenturer , uppbyggnad av nya nät och stöd till bestående nät .
Detta är bara några exempel .
Men det som är särskilt viktigt när det gäller Altener II-programmet är - anser jag - de nya åtgärderna för att underlätta att de förnybara energikällorna får genomslagskraft på marknaden , och de nya åtgärderna för att genomföra , åtfölja och övervaka gemenskapens strategi och gemenskapens åtgärdsplan .
Det föreligger nu ett arbetsdokument från kommissionens enhet rörande en kampanj för ett genombrott , vilken ju är en väsentlig beståndsdel i denna gemenskapsstrategi .
Det som här planeras är stöd på alla väsentliga områden i fråga om förnybara energikällor .
Detta Altener-program måste verkligen åtfölja och stödja denna kampanj .
De totala investeringskostnaderna för kampanjen har beräknats till ca 30 miljarder euro .
Därav skall 75 - 80 procent komma från privata källor , och härtill kommer allmänna medel från medlemsstater och regioner .
Här kan Altener-programmet ge viktiga nya impulser för investeringar , underlätta dem och hjälpa oss så att vi verkligen kan uppnå vårt mål beträffande miljöskydd , ekonomi och nya arbetstillfällen .
Herr talman , fru kommissionär !
Även jag vill tacka Langen för det goda arbete han lagt ned i detta viktiga ämne .
Det slutresultat av förlikningen avseende Altener-programmet som förlikningskommittén lagt fram är efter ett antal svåra turer åtminstone nöjaktigt .
Största delen av parlamentets ändringsförslag har beaktats , och som en positiv sak måste man konstatera att finansieringsbeloppet för programmet höjts till 77 miljoner euro .
När det gäller ökad användning av förnybara energikällor har unionen ambitiösa mål .
I förhållande till dessa mål är anslaget emellertid mycket litet .
Det måste användas till pilotprojekt , forskning , informationsutbyte samt till att bilda positiv opinion för användningen av förnybara energikällor .
Huvudansvaret för att öka användningen av förnybara energikällor vilar på medlemsstaternas axlar .
Förhoppningsvis väcker detta program medlemsstaterna till att bedriva en beslutsam verksamhet för att öka användningen av förnybara energikällor .
Men även unionen måste i framtiden öka sin egen satsning för att främja användningen av förnybara energikällor och se till att den förnybara energin utan hinder kan komma in på marknaden .
Att främja användningen av förnybara energikällor är särskilt viktigt med tanke på miljön .
Unionen kan inte uppnå sina miljömål om man inte aktivt ökar användningen av förnybara energikällor .
De förnybara energikällorna minskar beroendet av importerad energi och ökad användning av dem förbättrar konkurrenskraften .
Europa kan också uppnå en ledande position inom den industri som levererar de utrustningar som behövs för att använda förnybar energi .
Man måste också komma ihåg att användningen av förnybara energikällor har en positiv inverkan på den regionala utvecklingen och sysselsättningen .
Även jag vågar nämna torven .
Torven finns inte med på listan över förnybara energikällor .
Den är dock åtminstone i Finland en viktig , långsamt förnybar energikälla som används på ett hållbart sätt .
Jag hoppas att den i framtiden kan tas med på listan över förnybara energikällor .
Fru kommissionär , kära kolleger !
Gruppen De gröna gläds åt den överenskommelse som gjorts och vårt tack går till alla dem som förhandlat så bra för ett ändringsförslag som De gröna nästan var upphovsmän till .
Det är intressant för mig , som är ny här i parlamentet , att konstatera att man i budgeten planerar för hundratals miljoner euro per år för tobaksodling .
Det är en begränsad sektor av ekonomin som nästan inte skapar någon sysselsättning , som inte är konkurrenskraftig på världsnivå .
Jämfört med detta konstaterar jag de summor som står på spel för förnybar energi som inte bara är en ekologisk beståndsdel utan också är förutbestämd att få en avsevärd ekonomisk uppgång .
När man ser de marknadsandelar som små länder såsom Danmark lyckats förvärva på detta område , tack vare att de var de första på marknaden , tror jag det manar till eftertanke och att vi på lång sikt verkligen måste öka budgeten för förnybar energi .
Ett sista ord när det gäller programmet : Jag tror att det är mycket viktigt att de förnybara energikällorna , om de skall kunna utvecklas på lång sikt , är förankrade i regionerna där de kan bidra till ekonomin och till att skapa sysselsättning .
Om 50 procent eller mer av energimixen skall kunna komma från förnybara energikällor kan man inte nöja sig med vissa hot spots som på kort sikt blir mer lönsamma .
Herr talman !
Jag vill inleda med att gratulera herr Langen för hans arbete .
Aktiviteterna inom ramen för Altener-programmet kommer att främja förnybara energikällor och jag anser att sådana program förtjänar finansieringsstöd på utvecklingsstadiet då de erbjuder enorma kommersiella möjligheter i framtiden .
Av detta skäl är jag särskilt glad att se att pengarna satsats på små och medelstora företags projekt .
De internationellt överenskomna målen för minskade utsläpp kan inte uppnås genom dessa program enbart .
I detta hänseende måste man komma ihåg att energipolitiken förblir inom ramen för nationella befogenheter .
Det är ytterst viktigt att de nationella regeringarna ger sitt fulla stöd för att få en effektivare energianvändning och för att utveckla förnybara energikällor .
Jag är förtjust över att Irland nyligen meddelade att man där kommer att använda 125 miljoner irländska pund för att utveckla en miljömässigt hållbar energisektor .
Jag hoppas att Altener-programmet skall medverka och leda till fler initiativ .
Såsom korrekt fastslås i den slutgiltiga texten kan åtgärder som dessa spela en roll för att minska regionala skillnader .
Jag kan intyga att jag redan har mottagit bevis på stort intresse för Altener-programmet från min egen valkrets Leinster , en region som till en betydande del ligger inom Irlands enda mål 1-region .
Jag stöder alla insatser för att minska klyftan inom ekonomisk utveckling av infrastrukturbestämmelser , inklusive energisektorn .
Kort sagt , vi står inför en stor utmaning för att klara av våra åtaganden att begränsa utsläppen av växthusgaser från energisektorn enligt Kyoto-protokollet medan vi samtidigt främjar tillväxten i våra ekonomier .
Altener-programmet skall vara ett värdefullt bidrag till medlemsstaternas samlade insatser .
Herr talman , herr föredragande , kära kolleger !
Såsom vår föredragande erinrade om står vi nu vid slutet av en lång och svår förlikning med rådet om Altener-programmet .
Föredraganden erinrade om att det ekonomiska totalanslaget som rådet föreslagit ursprungligen var 74 miljoner francs medan kommissionen hade föreslagit 81,1 miljoner , ett belopp som Europaparlamentet stödde .
Ett första förlikningsmöte misslyckades , eftersom rådet då bara godtog en ökning på 1,9 miljoner euro .
Vi kunde inte godkänna ett sådant förslag som ifrågasatte Europaparlamentets befogenheter .
En andra förlikning gjorde det möjligt att öka på med 1,1 miljoner euro ytterligare för att uppnå denna kompromiss på 77 miljoner .
Trots en ökning på 3 miljoner i förhållande till det ursprungliga förslaget , beklagar jag personligen ännu en gång att de ekonomiska medlen inte är i nivå med de uttalade ambitionerna och att rådets strävan efter sparande i denna situation skiljer sig alltför mycket från dess uttalanden till förmån för säkerhet när det gäller energiförsörjning , skapande av sysselsättning samt miljöskydd som också är utmaningar som måste lösas .
Den förnybara energin utgör ett obestridligt medel för att uppnå dessa målsättningar .
Trots de förbehåll jag uttryckt om den svaga ekonomiska tilldelningen stöder jag ändå personligen kompromissen , på grund av programmets innehåll , ett innehåll som Europaparlamentet aktivt bidragit till eftersom detta område efter att Amsterdamfördraget trätt i kraft omfattas av medbeslutandet .
Man bör därför i stort sett med raden av genomförda och föreslagna åtgärder kunna närma sig målsättningen på 12 procent förnybar energi år 2010 , dvs. en fördubbling , om alla anslag , inklusive de statliga , följer med .
Detta program är tillsammans med programmet Save II , med införlivandet av miljödimensionen i energipolitiken , grunden för en verklig gemenskapsstrategi för att uppnå egen energi och samtidigt minska vårt beroende.Avslutningsvis , herr talman , tillåter jag mig också att betona att det utöver de åtgärder som föreslås också skall finnas lagstiftningsåtgärder och framför allt konsekventa budgetar för att åtfölja denna politiska vilja .
Och jag slutar naturligtvis med att lyckönska herr Langen , vår föredragande , för hans arbete , liksom samtliga medlemmar i utskottet och förlikningskommittén . - Herr talman , mina damer och herrar !
Jag vill börja med att uttrycka min glädje över den överenskommelse som har uppnåtts angående programmet Altener II i förlikningskommittén och ansluta mig till de uttalanden som har gjorts av tidigare talare , och givetvis påpeka att denna överenskommelse kommer att innebära att programmet Altener inom kort tas med i ramprogrammet för energi .
Allt detta kommer att leda till en ökad samordning , insyn och effektivitet i våra energiprogram , i vilka även programmet Save måste införlivas , vilket vi snart kommer att diskutera .
Jag anser att parlamentets arbeten under den här perioden har hållit hög standard , och därför gratulerar jag föredragande Langen och även de olika talare som har hållit anföranden , både i kommissionen och här i parlamentet .
Det är uppenbart att det har förts diskussioner , vi blev tvungna att söka förlikning , precis som föredraganden och Caudron påpekade för en stund sedan , för under det första mötet uppnåddes inga resultat , och man blev därför tvungen att samlas en andra gång , trots att siffrorna inte heller var överdrivet höga .
Men jag anser att vi till slut lyckades uppnå ett rimligt avtal som i likhet med alla avtal inte är fulländat , men som jag tror gör det möjligt att fortsätta med de projekt som vi hade på gång .
Därför vill jag upprepa mina gratulationer till föredraganden Langen för det arbete han har utfört , tacka alla talare och naturligtvis lovorda vice ordförande Provans agerande under förlikningsförfarandet som i stor mån bidrog till att uppnå ett positivt resultat .
Jag vill även lovorda rådets förnuftiga och flexibla attityd .
 
Save Nästa punkt på föredragningslistan är betänkande ( A5-0010 / 2000 ) av Ahern för Europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets beslut om att anta ett flerårigt program för att främja en effektiv energianvändning - Save ( C5-0334 / 1999 - 1997 / 0371 ( COD ) ) . . - ( EN ) Fru talman !
Jag vill tacka rådet och kommissionen för ett bra och omsorgsfullt förlikningsförfarande där alla var vid gott humör vilket inte alltid är fallet .
Det är ett nöje för mig att säga att jag anser slutresultatet av förlikningen som mycket tillfredsställande för parlamentet då den gemensamma texten innehöll alla dess ändringsförslag antingen hela texten eller i omformulerad form .
Det belopp som slutligen anslogs till programmet är också en betydande förbättring mot rådets förslag vid den andra behandlingen som vi ansåg som helt oacceptabelt och vi har lyckats få betydande framgång där .
Jag föreslår därför att denna kammare antar förslagen för Save-programmet och slutsatsen vid förlikningen vid tredje behandlingen .
Jag vill påminna kammaren om att vid andra behandlingen godkände parlamentet detta betänkande innehållande åtta ändringsförslag , inklusive ett återinförande av kommissionens ursprungliga budget .
Kommissionen godkände fem av de föreslagna ändringsförslagen , inklusive budgetanslaget , och jag tackar kommissionen för deras fortsatta stöd om budgeten under förlikningsförfarandet då det som rådet hade föreslagit var oacceptabelt .
Under förfarandet kom man överens om vilka undersökningar och insatser som skulle planeras , genomföras , kompletteras och utvärdera gemenskapsinsatserna .
Kompromissformuleringar enades man om för fem andra ändringsförslag inklusive lagstiftnings- och icke lagstiftningsåtgärder och inrättandet av lokala energicentra och , något mycket viktigt , energikontrollsystem en som skall följa upp utvecklingen av ökad energieffektivitet .
Jag hoppas att ni alla skall hålla med om att detta är en viktig utveckling .
Frågan om det finansiella anslaget försvarades hårdnackat av parlamentet ställt mot rådets mycket låga öppningserbjudande .
I varje fall fick vi lova att hålla flera sammanträden innan rådet slutligen höjde beloppet avsevärt .
Vi fick en ökning med 2 miljoner mot deras första förslag , vilket var en betydande höjning som jag kan rekommendera er och som kommissionen bekräftade skulle räcka för att den skulle kunna genomföra programmen .
Detta var ett viktigt ställningstagande för oss .
Jag skulle dock vilja framföra att det är och har alltid varit en mycket blygsam budget och därför är finansieringen för detta program mer symbolisk än reell .
Finansieringen för att spara energi görs fortfarande huvudsakligen av medlemsstaterna .
Vi måste komma ihåg det när vi godkänner detta program .
Om det är fråga om mer symbolism än realitet i fråga om det som vi kan uppnå på gemenskapsnivå är det synd för det finns mycket entusiasm på lokal nivå för åtgärder , däribland gemenskapsåtgärder , för energibesparing .
Ett område där gemenskapen kan hjälpa till är att skapa kontakter mellan lokala aktörer så att de inte behöver starta om från början i varje region .
Vi har en betydelsefull roll att spela i gemenskapen inom Europeiska unionen i detta avseende .
Save är det enda program som täcker hela gemenskapen och som är avsett att främja en rationell energianvändning .
Det är inriktat på icke tekniska områden för att skapa energieffektiva infrastrukturer och ändamålet med programmet är att skapa en miljö för att främja investeringar och en effektiv energianvändning .
Här behöver vi inse att det även finns en marknadsmöjlighet inom industrin för energibesparingar .
Vi har hört en massa om konkurrenssvårigheter inom förnybara energikällor men energieffektivitet sparar pengar för företag , sparar pengar överallt i själva verket , och därför bör det inte finnas problem här .
Det är något som vi alla kan stödja .
Jag måste säga , liksom moderskap , även om vi alla stöder det , gör vi ibland mycket lite i det stora hela och rent konkret för att hjälpa mödrar eller människor som är intresserade av energibesparing .
Vi kan göra ganska mycket mer med hänsyn till att vi har gjort stora åtaganden för att minska utsläppen av koldioxid och växthusgaser och för att minska beroendet av energiimport .
Vi vidtar inte de åtgärder som medborgarna önskar .
Vi visar inte på sambandet så att medborgarna verkligen kan göra något konkret i hemmet eller på sina kontor eller i industrin för att stödja åtgärderna mot globala klimatförändringar .
Om vi kan föra fram detta budskap skulle det vara en mycket intressant sak att göra .
Jag vill återigen tacka alla som hjälpte till i detta förlikningsförfarande . - Fru talman , mina damer och herrar !
Jag vill åter igen tacka fru Ahern för hennes arbete som föredragande av detta förslag , för hon har i samarbete med övriga parlamentariker bidragit till att man slutligen uppnått ett högst rimligt resultat , som i vissa avseenden även förbättrar en del av kommissionens förslag och naturligtvis det som rådet till en början hade godkänt ur budgetsynpunkt .
Precis som Ahern så riktigt sade är både budgeten för Save- programmet och den för Altener-programmet , i första hand symboliska budgetar , för den tyngsta bördan bär länderna , unionens stater , regionerna och även i vissa fall kommunerna .
Hur som helst innebär inte dess begränsade volym att den upphör att ha det viktiga symboliska värde som förutsätts av det faktum att det inom gemenskapen som helhet finns en vilja att stödja denna typ av åtgärder som bidrar till att vi verkligen uppfyller våra löften från Kyoto och dessutom till att vi uppnår ett större mångfald i våra energikällor , en ökad säkerhet i vår energiförsörjning och , som i fallet med Save , att vi närmar oss en lägre konsumtion , ett mer effektivt utnyttjande av energin , och därigenom bidrar till att nå de uppsatta målen .
Dessutom står vi nu i samband med dessa program , det vill säga Save-programmet för en effektiv energianvändning och Altener-programmet för förnybara energikällor , inför en mycket viktig teknisk utmaning , som ur ekonomisk synvinkel kan komma att innebära stora möjligheter för industrin och även för skapandet av sysselsättning i våra länder , och därigenom i hela unionen .
Vad beträffar den parlamentariska behandlingen , vill jag upprepa mitt tack till alla de som har agerat och talat , och huvudsakligen föredraganden , för i det förslag som har godkänts av rådet har de flesta av parlamentets ändringsförslag tagits med , praktiskt taget samtliga i det här fallet , om än med vissa ändringar , och jag vill tacka för att man dessutom har lyckats förbättra det första erbjudandet vad medlen beträffar .
Det har man lyckats göra med hjälp av nya pengar , så som vi den gången sade , och man har lyckats göra det och samtidigt bevara parlamentets förmåner och behörighet .
Från kommissionens sida sett , i detta spel institutionerna emellan , anser jag att det är viktigt , och jag har nöjet att få poängtera detta .
Jag vill upprepa mitt tack till alla som har talat , i synnerhet till vice ordförande Provan , för hans föredömliga agerande under denna debatt , framför allt under förlikningsprocessen , till ordföranden i utskottet för industrifrågor , utrikeshandel , forskning och energi , och även till föredragande Ahern , samt till alla de ledamöter som har deltagit i arbetet .
Tack , fru kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11 .
 
Kultur 2000 Nästa punkt på föredragningslistan är betänkande ( A5-0009 / 2000 ) av Graça Moura för Europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets beslut om att inrätta ett enhetligt instrument för finansiering och programplanering för kulturellt samarbete ( Kultur 2000-programmet ) C5-0327 / 1999 - 1998 / 0169 ( COD ) ) .
Fru talman !
Trots artikel 151 i Amsterdamfördraget har kulturen varit den sektor som dragit det kortaste strået i den krympande programapparaten och när det gäller de finansiella , tekniska och mänskliga resurser som mobiliserats för det europeiska projektet .
Man kan säga att de mål som för 50 år sedan var grundvalen för det " europeiska hus " vi i dag lever i var mera specifikt ekonomiska och sociala .
Man kan också säga att den europeiska politiken under de här fem årtiondena har påverkats av många olika impulser i de mest varierande konjunkturer och av många olika skäl .
I sinnet hos Europas grundare måste det dock ha funnits en civilisationstanke som fick oss att vilja skapa hållbara förutsättningar för fred .
En sådan tanke är baserad på omfattande kulturell mångfald .
Ett Europa med en nationell identitet kan leva i fred och välmåga under väldigt lång tid , en förutsättning är dock att vitaliteten i den kulturella mångfalden bevaras , att den förbittrade småaktighet och agressivitet som i regel leder till överdriven nationalism elimineras .
För att möjliggöra detta är det absolut nödvändigt att vi har kunskap om varandra och att vi utgår från värden av sann mänsklighet och tolerans när det gäller de artistiska och kulturella uttrycken , uttryck som slår rot i den bördiga europeiska myllan och som talar om vad som är det mest storsinta och sinnrika i den mänskliga själen .
För att denna vetskap och denna utgångspunkt fullt ut skall bli möjlig måste vi följaktligen enas om hur kulturen i den europeiska demokratin skall uppfattas .
Den faktiska konvergensen , den ekonomiska och sociala sammanhållningen , kampen mot arbetslöshet och utanförskap och till och med konkurrensen är tvivelsutan förutsättningarna för att skapa större jämlikhet , större tillväxt , bättre livskvalitet och bättre möjligheter för de europeiska medborgarna .
Den gemensamma försvars- och säkerhetspolitiken kan säkert också förstärka den europeiska identiteten och bekräftelsen i världen .
Den politik som bedrivs för värnandet om de mänskliga rättigheterna är också tvivelsutan ett universellt projekt .
Kan man inte i det kulturpolitiska arbetet ge allt detta en djupare mening och klarare kriterium , så kan varken Europa eller den europeiska demokratin gå mycket längre .
Det är genom kulturen och bara genom den som miljontals medborgare kan känna sig som européer och odla , bearbeta och fördjupa känslan av att tillhöra Europa .
Fru talman , det är detta vingslag som har saknats i den europeiska politiken .
Man talar om kultur , om kulturellt samarbete , emblematiska åtgärder , stora initiativ , nätverk av agenter och kulturella operatörer , men man undviker noggrant att hänvisa till den kulturella politiken vid de europeiska institutionerna , som för övrigt inte på något sätt skulle kollidera med subsidiaritetsprincipen .
Samtidigt talar man , ibland retoriskt uttrycksfullt , om kulturens betydelse för det europeiska projektet , men löjliga summor reserveras för program som beständigt och regelbundet borde betjäna mer än 300 miljoner människor och ge dem tillträde till ett fädernearv som tillhör dem och som skulle kunna väcka en aktiv och interaktiv lust för de stora värdena och de stora skapelserna .
Europas medborgare , som vi här företräder , har rätt att av unionens institutioner kräva en fastare , effektivare och mera europeisk hållning .
Sådana överväganden kan ses som en början till kammarens erkännande av det gemensamma projektet Kultur 2000-programmet , godkänt av förlikningskommittén den 9 december .
Kom ihåg att Kultur 2000 ger oss ett unikt finansierings- och programplaneringsinstrument för det kulturella samarbetet .
Resultatet av förlikningen var tillfredsställande när det gäller nästan alla de ändringsförslag som godkändes vid andra behandlingen , den grundläggande förståelsen hos parlamentet kan därmed skäligen anses rättfärdigad , särskilt beträffande den politiska prioriteringen att skapa förutsättningar för att åtgärderna i Kultur 2000 skall nå så många medborgare som möjligt .
Beträffande budgetaspekterna så mötte parlamentets delegation rådets okuvlighet när det gäller den anslagsökning på 167 miljoner euro som man till en början hade förutspått .
Man stannade vid en från den här ståndpunkten sett förmildrande lösning , för övrigt genomförbar enbart tack vare kommissionär Viviane Redings försök att finna en konstruktiv lösning .
Kommissionen kunde därmed förbinda sig att före den 30 juni 2002 lägga fram ett betänkande om programmets funktion där man uttalar sig om de tillgängliga finansiella resurserna i fråga om kapacitet eller inkapacitet och där man föreslår en eventuell revidering av den punkten .
Vi får dock inte dölja att framgången av ett sådant förslag i korthet beror på om man under tiden har funnit någon institutionell mekanism som motsvarar den egentliga meningen med termen " förlikning " .
Avslutningsvis uppmanar jag kammaren att ge det gemensamma av förlikningskommittén godkända projektet Kultur 2000-programmet sitt absoluta stöd och jag önskar programmet all välgång .
Fru talman !
Jag tror egentligen att vi inte hade behövt tala mer om det , ty vi har redan sagt allting under den senaste debatten .
Tyvärr har ju ingenting ändrats i fråga om det faktum att rådet alltid talar om kultur , men inte ger ut några pengar för kultur .
Vi har en känsla av , och är egentligen övertygade om , att medlemsstaterna skulle uppskatta om de kunde stryka det som de 1992 skrev in i Maastrichtfördraget .
Ty ingen vill egentligen verkligen ge ut pengar för kultur .
Tyvärr är det så .
Det måste vi konstatera .
Jag vill tacka föredraganden , som verkligen oförtröttat har arbetat med detta omfattande ärende , naturligtvis i samarbete med kommissionären .
Vi måste nog notera att vi egentligen har uppnått vårt mål beträffande innehållet , men naturligtvis inte beträffande finanserna .
I en sådan förlikning , där man å ena sidan verkligen måste uppnå enhällighet , känner man sig maktlös .
Det är egentligen inte någon rättvis basar !
Det finns alltid människor där som kan avvisa allting , och å andra sidan står vi och tigger om lite mer för kulturen .
Det är egentligen vanhedrande , det som vi gör där !
Det är en förskräcklig arabisk basar , med ojämna förutsättningar .
Det gläder oss ändå att detta program har blivit sådant som vi önskade .
Det motsvarar det som medborgarna förväntar sig av oss .
Vi stöder små och medelstora arrangemang , inte de stora arrangemangen , vi gör tillgången till det enklare för den enskilde medborgaren och även de mindre aktörerna ; jag tror att det faktum att kulturen i dag ju tillsammans med utbildning och ungdom befinner sig i en kommissionärs hand , också borgar för att det skapas mer synergi mellan dessa tre program , som ju är utpräglade program för medborgarna i Europeiska unionen .
Om man tar alla pengar och åstadkommer synergieffekter , då kan man var litet tillfreds , men också bara litet grand .
Jag önskar att vi med dessa mindre summor uppnår många effekter .
Fru talman !
Jag håller med om de stora ord som fick inleda föredragandens anförande , men jag måste få tillägga att jag under förlikningen har blivit lite besviken på rådet .
Å ena sidan vägrade man fortfarande att acceptera begreppet " europeisk kulturpolitik " och liknande begrepp , bland annat genom att förringa det som står i fördragen , och man har endast definierat begreppet " kultur 2000 " som ett instrument för ett kulturellt samarbete , och mer än så blir det inte .
Å andra sidan har man visat sig helt omedgörlig beträffande den finansiering som parlamentet har begärt , som gällde en minimifinansiering .
Nåja , det vore orättvist att påstå att det sista rörde rådets fjorton medlemmar , för det var bara en , Nederländerna , som i första hand visade sig omedgörlig .
Det har än en gång visat sig att en förlikning är oförenlig med kravet på enhällighet i rådet .
Ett sådant krav gör i princip en förlikning omöjlig och inverkar dessutom på den parlamentariska institutionens värdighet .
Fru talman , dessa överväganden får emellertid inte dölja det faktum att denna text som i sin helhet kommer att bli föremål för omröstning i morgon , och som vi socialister kommer att rösta för , kommer att innebära igångsättandet av ett av Europeiska unionens viktigaste program .
Genom att agera på det kulturella området , skapar vi Europas själ , inte minst i det här fallet med de fantastiska gemenskapsprogram som utgör " Kultur 2000 " .
De senaste åren har dessa blivit de mest accepterade programmen bland de mest dynamiska och yngsta medborgarna i Europeiska unionen .
Slutligen vill jag nämna det starka intryck som föredragande Graca Moura som individ har gjort på mig : hans kunskap , hans eftertanke , hans intellektuella nivå visar , anser jag , att han är den bästa föredraganden som detta betänkande hade kunnat få .
Gratulerar !
Till sist vill jag gratulera kommissionär Reding , vice talman Imbeni samt Gargani , ordförande i utskottet för kultur , ungdomsfrågor , utbildning , medier och idrott , för den bestämda och kloka hållning som de , var och en i sin roll , har intagit under hela förlikningsprocessen .
Fru talman , fru kommissionär , herr föredragande !
Jag skulle vilja börja med att tacka Graça Moura så hjärtligt för hans fantastiska insats under behandlingen av programmet Kultur 2000 .
Det har redan sagts och vi har diskuterat det flera gånger , kultur är naturligtvis otroligt viktigt som ett självständigt område , det vill jag betona igen , men också som ett utmärkt instrument för att vidarebefordra den europeiska tanken och kulturen är mycket viktig för medborgarna .
Det får vi absolut inte glömma bort .
Det europeiska stimulans som ges ut genom det här programmet medför otroligt mycket , särskilt för små språkområden som t.ex.
Nederländerna där det inte endast gäller nationella möjligheter men de behöver också stödjas , framförallt genom språket .
I dag har vi kommit fram till slutet av en lång resa .
Jag skulle ändå helt kort vilja , precis som andra gjort , gå in på det otydliga och främst ovälkomna förfarandet .
Medbeslutande och enhällighet är som en orm som biter sig själv i svansen .
Det finns inte mycket att förhandla om i fall en av parterna på förhand säger : vi kan prata om allt men budgeten står fast .
Nu har , och det vill jag ändå också säga när det gäller Nederländerna , förhandlingarna om det redan ägt rum i ett tidigare skede .
Resultatet är 30 procents tillväxt , så vi är inte helt olyckliga över resultatet .
Det är naturligtvis alltid bättre , och det skall jag alltid yrka för , att anslå mer pengar och även något snabbare .
Ändå så tror jag att det här programmet erbjuder goda chanser för flera olika program .
Jag skulle vilja betona att kultur inte enbart får stöd från den här fonden .
Kultur består inte enbart av kultur utan även av många andra områden .
I strukturfonderna finns också mycket pengar tillgängliga för kultur och det måste vi ju också ta i gott beaktande .
Lyckligtvis är jag ledamot i utskottet för regionalpolitik .
Jag skall alltså själv se till att det också sker i stor utsträckning .
Jag tror att vi även tagit ställning för att instämma i att budgeten är tillräckligt omfattande , om det inte går igenom så är det ju ändå dåligt för medborgaren .
I det avseendet har jag också alltid stöttat föredraganden .
Jag tycker dock att det , och det säger han också alltid , vid den kommande regeringskonferensen behöver göras en ändring i medbeslutandeförfarandet , då behövs ingen enhällighet .
Vi är mycket positiva över de många förbättringar som skett .
Inga megaprojekt längre , utrymme för kulturella nätverk , god uppmärksamhet för läsfrämjande åtgärder , översättning , översättarhus , mycket viktigt för de mindre språkområdena .
Jag vill verkligen lyckönska föredraganden och även Reding till Kultur 2000 .
Det enda som återstår för mig att säga är : nu sätter vi igång .
Fru talman !
De kolleger som har talat före mig har sagt det mesta , och jag tror att det finns en samstämmighet bland grupperna i Europaparlamentet liksom bland alla oss i utskottet för kultur , ungdomsfrågor , utbildning , medier och idrott .
Även jag skall säga att det är med ett mycket tungt hjärta som jag kommer att rösta för detta gemensamma förslag till rådets och Europaparlamentets beslut .
Inte på grund av att våra företrädare , vår föredragande och ordföranden Gargani , inte har uträttat ett enastående arbete - det har lagt ned enormt mycket arbete - , inte på grund av att jag har några stora invändningar mot den ståndpunkt som kommissionär Reding har vidhållit - jag tycker att hon inom de ramar som hon hade vidhöll en mycket positiv ståndpunkt - , utan på grund av rådets negativa och oacceptabla inställning .
Det är en skam !
Denna siffra , 167 miljoner euro för så många år , är en skam för Europeiska unionen !
När vi bokstavligen tvingas att kväva teatergrupper , unga musiker , innovativa verksamheter inom konst och litteratur , att kväva dem och hålla god min och ge femtioelva avslag , med resultatet att de uppfattar Europa som någonting främmande , någonting motsträvigt , någonting negativt och någonting fientligt i sina ansträngningar att skapa kultur , ansträngningar som Europeiska unionen måste stödja - för vår väg är inte bara euron , inte heller bara utvidgningen eller egoistiska geostrategiska hänsyn ; den är att ge en kulturell blomstring till den europeisk integrering - , är denna utgång beklaglig .
Och så länge som vi har kvar enhälligheten och så länge som en regering , som Nederländernas regering i går , kan fastställa de där 167 miljonerna med ett ultimatum och så länge som en regering med Haider i övermorgon kan tala om för oss vilka kulturella verksamheter vi skall ägna oss åt , kommer vi inte att komma framåt .
Därför är det mycket viktigt för regeringskonferensen att det fattas viktiga beslut och att det kommer till stånd en ändring , så att Europaparlamentets ansträngningar att få till stånd en viktig kulturell blomstring inom det europeiska området befrias från enskilda regeringarnas tvångströjor .
Fru talman !
Jag delar helt de värderingar som har framförts av föredraganden och jag vill också tacka ordföranden för utskottet för kultur , Gargani , för det berömvärda arbete han utfört under en medlingsprocess som även varit ganska komplicerad .
Utan tvekan finns det behov av att förenkla och förstärka tidigare program men alla hoppades att programmet Kultur 2000 skulle kunna bidra till att till exempel främja varje kultursektors särart , och även - eller framför allt , bör man kanske säga - de sektorer som inte är så kända .
Vi hoppas att detta skall inträffa , åtminstone när det gäller finansieringen .
Vi tror mycket på värdet av kulturella handlingar , även när det gäller bidragen till ett folks sociala och ekonomiska tillväxt .
Och Europa kan fullt ut konkurrera med resten av världen genom att till fullo återupptäcka sina rötter , genom att förverkliga det gemensamma kulturella nätverket , genom att utnyttja och återge värdigheten åt de kulturella och språkliga öar som hittills varit mindre kända .
När det gäller den stora pedagogiska uppgift som Europeiska unionen står inför i samband med den kulturella dimensionen , är finansieringen en av de tydligaste begränsningarna när det gäller programmet - det har vi fått höra flera gånger - och något som pekar på att man inte har helt förstått - åtminstone gäller det rådet , men sannerligen inte kommissionären - betydelsen av denna kulturella uppgift : detta visar även dokumentet som prioriterar de ekonomiska faktorerna framför den sociala integrationen .
En allsidig tillväxt av Europeiska unionen och medvetenhet om vad det innebär att vara europeiska medborgare : det är därför vi anser att projektet Kultur 2000 , även när det gäller finansieringen , skulle kunna lämna viktiga bidrag till detta stora gemensamma mål .
Fru talman !
Jag vill öka kvällens enhällighet och säga att jag stöder godkännandet av Kultur 2000 och framför mina tack till föredragande , Graca Moura , som efterträdde vår förra kollega Nana Mouskouri .
Båda har gjort ett förstklassigt arbete .
Vid sidan av den debatt vi hade tidigare i dag kanske kultur inte verkar vara så viktig men den är det och vi måste vara varsamma i Europaparlamentet så att brådskande frågor inte går före vad som är viktigt .
Varför anser jag att kultur är viktig ?
Jo , i enkla ekonomiska termer främjar europeisk kultur verkligt välstånd .
Var skulle Europas turistindustri befinna sig utan rikedomen i vår kultur ?
Men viktigare än det , kulturaktiviteter är det som gör människosläktet civiliserat .
Kulturen är grunden för vår tro på demokrati och ett icke kulturellt samhälle kan inte upprätthålla tolerans och frihet och demokrati .
Kulturell mångfald är viktig och den är hotad .
Men hotet kommer inte från Europa .
Många människor i mitt land säger att de uppfattar att brittisk kultur hotas exempelvis från Portugal , Tyskland , Finland , för guds skull .
Vi dricker ju portvin och vi tycker om tyskt öl och vi använder till och med finsk bastu men det är inte från Europa som kulturen hotas .
Vad jag verkligen ser i hela Europa är folk som dricker Coca Cola , som äter hamburgare , bär baseballmössor , tittar på Hollywoodfilmer och ofta gör allt detta samtidigt .
Jag tror inte att protektionism och reglering är rätt metod för att försvara Europas kultur , men jag tror att vi ska ge en hjälpande hand när vi har möjlighet .
Det är vad Kultur 2000 handlar om .
Så jag säger till ministerrådet : Utvärdera verkligen ständigt detta program .
Gör vi tillräckligt mycket ?
Och jag säger till fru Reding , tack för det stöd och den hjälp ni har gett hittills , fortsätt göra ett bra jobb , vi står på er sida .
Fru talman !
Även jag vill varmt tacka föredraganden Graça Moura och kommissionsledamoten Reding för deras ansträngningar för att åstadkomma detta program .
Kultur 2000-programmet fick ju sin slutgiltiga form i slutet av förra året genom förlikningen mellan parlamentet och rådet .
Slutresultatet kan anses vara rimligt med tanke på att det krävdes ett enhälligt beslut i rådet för att godkänna programmet .
Det är önskvärt att man vid den kommande regeringskonferensen kommer fram till att införa beslut med kvalificerad majoritet även inom kulturens område .
Det är verkligen besynnerligt att lagstiftning där man tillämpar medbeslutandeförfarandet förutsätter enhällighet i rådet .
Det kulturella ramprogrammet ersätter de nuvarande programmen Kalejdoskop , Ariane och Rafael .
När man börjar genomföra programmet hoppas jag speciellt att möjligheterna för litteraturen och översättningen av böcker kan utnyttjas fullt ut .
Jag tror och hoppas att litteraturen bibehåller sin ställning trots den nya teknikens framfart .
Vi behöver den fördjupning som litteraturen erbjuder mitt i all kortsiktighet och ytlighet .
Litteraturen har likaså en stor betydelse när det gäller att förmedla vårt kulturarv , att öka kännedomen om varandra samt att omhulda den språkliga rikedomen och mångfalden .
I detta sammanhang är det speciellt angenämt att konstatera att EU : s ordförandeland strax efter att Sokrates- och Kultur 2000-programmet startats kommer att anordna ett möte där man skall dryfta bibliotekens ställning .
Jag hoppas att detta möte också skall uppmuntra kommissionen till att på ett aktivt sätt beakta biblioteken i informationssamhällets femte ramprogram .
Fru talman , fru kommissionär , herr föredragande , mina damer och herrar !
Någonstans sluts kretsen med dagens föredragningslista .
Vi har i dag talat mycket om Europa som en värdegemenskap , om tolerans , mänsklig värdighet , mänskliga rättigheter , ett positivt förhållande till utvidgningsprocessen , öppenhet och respekt för varandra .
Ungdoms- , utbildnings- och kulturpolitik är viktiga verktyg när man skall skapa dessa värden , skapa förtroende hos medborgarna i Europeiska unionen och skapa trovärdighet för Europeiska unionen gentemot medborgarna .
De finansiella medel som av rådet medgivits för kulturprogrammet står i ett slående motsatsförhållande till betydelsen av kultur- och utbildningspolitiken samt detta program för Europeiska unionens mål .
Kulturell verksamhet skapar identitet .
Kulturell verksamhet är ett uttryck för individualitet och den egna personligheten , den skapar kontakt och kommunicerar .
Vi vill ha ett brokigt Europa .
Vi vill ha ett Europa enligt principen mångfald inom enheten .
Vi vill att människorna skall lära sig förstå och uppskatta skillnaderna .
Av den anledningen har vi uttalat oss för en uppdelning av budgeten respektive anslag till de olika typerna av åtgärder .
Av den anledningen har vi avvisat den starka koncentrationen till stora nätverk och nätstrukturer , eftersom vi vill främja de små och medelstora enheterna , den individuella verksamheten , eftersom vi vill låta tusen blommor blomma .
Jag vill stödja de föregående talarna .
Det är en motsägelse - enhällighetsprincip , medbeslutandeförfarande och förlikningskommitté - om vi vill stärka kulturpolitikens principer för ett europeiskt medvetande och inte vill fortsätta att försvaga dem .
Fru talman , mina damer och herrar !
Som vi har hört , har alla våra grupper en gemensam politisk fiende , och det är rådet .
Utskottets för kultur beslut hamnar ju inte av en tillfällighet alltid i ett förlikningsförfarande , ty det är alltid något medlemsland i rådet som tar kulturen till gisslan för andra intressen .
Så visar sig enhällighetsprincipen vara ett första klassens blockadinstrument .
I nästan två år har man brottats för att uppnå en genomförbar kompromiss , innan Europaparlamentet nu äntligen kan ge grönt ljus .
Inte ens det faktum att de föregående programmen Kaleidoskop , Ariane och Rafael löpte ut kunde beveka rådet .
Det krävdes ett pilotprogram för att överbrygga detta .
Det har än en gång tydliggjort svagheterna i Europeiska unionens kulturpolitiska åtgärder .
Den politiska kampen om anslagsfördelningen och programutformningen står inte i någon proportion till volymen på stöden .
Av 410 framställningar år 1999 kunde bara 55 projekt med en mager totalvolym om 6,07 miljoner euro beaktas .
Beträffande föreliggande program var rådet inte berett att komma parlamentet till mötes med en enda euro !
Alltså stannar vi kvar på blygsamma 167 miljoner till år 2004 .
Det motsvarar utgifterna för ett enda medelstort tyskt operahus under samma period , medan denna summa här i Europa är avsedd för 29 länder i över 5 år .
Det är ett krasst missförhållande !
Alltså måste vi då vredgat finna oss till rätta med att vi åtminstone i fråga om innehållet har fått igenom en del .
Det har ju också redan lyckligtvis skildrats .
Hoppet kvarstår att det en dag kommer att bli möjligt att förmå rådet att ändra inställning .
Kanske kommer man ju också att begripa att Europeiska unionens kulturella aktiviteter inte utgör någon fara , utan en möjlighet !
Kulturellt samarbete - även detta har skildrats - bidrar sannerligen till att ge en identitet , mycket mer än alla viktiga transportdirektiv .
Att man främjar kulturen bemöts med allmän acceptans , vilket man sannerligen inte kan påstå om alla politiska beslut .
Vad är det alltså , frågar jag er , som rådet är ängsligt för ?
Fru talman !
Den som , i likhet med mig , har äran att vara ordförande för kulturutskottet kan inte annat än instämma i det som har sagts av diverse kolleger och jag kan inte låta bli att gratulera föredraganden och kommissionären , fru Reding , med vilken föredraganden har arbetet och som , även i förlikningen , har haft svåra stunder , har kämpat mot rådet , det har vi fått höra av alla .
Jag har kunnat konstatera hur starkt man har bekräftat principen om kulturens nödvändighet när det gäller det europeiska konstruktionsarbetet men med små möjligheter att tillfredsställa alla de krav som kommer från Europas olika stater .
Låt mig bara understryka mitt personliga beklagande över att man i slutändan inte har lyckats godkänna en revideringsklausul .
Vi har , det är sant , fru Redings villighet och långsiktiga mål , Reding som har engagerat sig personligen för att ta upp frågan på nytt , för att göra en heltäckande utvärdering om något år , och därmed få till stånd en ny situation .
De olika kulturprogram - Kaleidoskop , Ariane , Rafael - som har startats under de år som gått ersätts nu av ett enda program , Kultur 2000 , där - detta vill jag gärna understryka - föredraganden stigmatiserat en åsikt som borde få Europaparlamentet att tänka efter - vilket någon redan påpekat under eftermiddagen i dag - men som alltid understryker den stora betydelsen av att vara del av en stor gemenskap där kulturen är ett demokratiskt fenomen .
Detta är ingen tom retorik , utan snarare en ny typ av liberalism som förenar de europeiska staterna och som är en utmaning för Europaparlamentet och kommissionen .
Vi har enats i den här frågan och det resultat som vi i dag har uppnått , trots den bristfälliga finansieringen , tror jag kan göra så att denna strategi och denna möjlighet för Europa verkligen får en bred lansering , en strategi som kommer att bli avgörande för såväl ekonomin som utvecklingen : med andra ord kulturen , ett institutionellt och organisatoriskt faktum som en förutsättning för den ekonomiska utvecklingen , och inte tvärtom , som Europa av tradition tyvärr har haft för ovana att se det under de år som gått .
I första hand handlar det om människan , i första hand handlar det om kulturen , och den kulturen kan avgöra den ekonomiska utvecklingen .
Låt oss begrunda detta resultat , låt oss vara glada och låt oss ge oss själva stor frihet att utforma en användbar strategi .
Fru talman !
Får jag först och främst tacka herr Graça Moura för att ha vävt sin väg genom de ganska hårda vävnader och trådar som denna förlikningsvävnad bestod av .
Det förefaller mig när vi inledde förliknings- förfarandet för Kultur 2000 att det är helt passande att ha en poet att leda oss i vår strävan .
Då dessa förlikningar inte utvecklas i helt rak kurs måste vi på nytt tacka vice talman Imbeni för hans föredömliga förhandlingsskicklighet på det invecklade området för att se till att kulturanslag sprids ut på ett klokt sätt och ges till oss i vår gemenskap .
Jag tycker att den huvudfråga som detta parlament , kommissionen och rådet står inför verkar vara : Vad är Europa ?
Vad betyder Europa och vad ger Europa oss utöver parametrarna för våra nationella gränser ?
Europa är dess folk , dess historia och nu dess gemenskap .
Skälet till varför Kultur 2000 är så viktig för oss är emellertid detta : Jag skall slå vad om det när vi ställer frågan - ' Vad är Europa ?
Vi svarar med att säga : " Det är vår konst , det är vår litteratur och det är vårt arv . "
Det är vad Kultur 2000 står för .
Detta program står för möjligheten att bibehålla en europeisk identitet på 2000-talet , en identitet som saknar ekon av splittring , av krig , av fattigdom , av möjligheter , av fattigdom i verkligheten .
Och mer än detta - och detta är mer vardagligt , fru talman , innebär det att vi har förmåga att lära från tidigare politiska initiativ genom att tillämpa dem i nya program som är innehållsrika , som täcker flera områden och som är till nytta för våra kreativa industrier i den utsträckning som de nu behöver .
Det främjar rörlighet och öppnar dörrar till kultur för de socialt missgynnade och utslagna .
Det enda jag beklagar är att vi inte har tillräckligt med pengar för att stödja detta program i överensstämmelse med våra förhoppningar och så att vi kan säkerställa att vi kommer att kunna nå ända fram . .
( FR ) Fru talman , mina damer och herrar !
Vi har nu kommit till slutet på en lång väg .
Efter förlikningsetappen kan våra institutioner numera formellt anta det nya ramprogrammet " Kultur 2000 " .
Vi förfogar då över ett instrument som gör det fullständigt möjligt att under de fem kommande åren utveckla en tydlig och väl strukturerad och , det är jag säger på , lönsam åtgärd , till förmån för kultursektorn .
Det är med tillfredsställelse jag i dag här välkomnar denna happy end och jag tackar er .
Jag tackar alla dem som här i parlamentet arbetat för att en bra avslutning på förlikningen kunnat bli möjlig .
Jag vill uttrycka mitt tack särskilt till utskottet för kultur , ungdomsfrågor , utbildning , medier och idrott och bl.a. dess föredragande Graça Moura , dess ordförande Gargani , till Europaparlamentets delegation och de ansvariga för de politiska grupperna , till förlikningskommittén och dess ordförande Imbeni .
Alla har bidragit konstruktivt , rättvist och beslutsamt .
Under hela denna förhandling har de varit till stor hjälp och det måste sägas att den svåra , ibland smärtsamma , förhandlingen ändå genomförts på rekordtid .
Vi har nu ett ramprogram , det första i detta slag för kultursektorn , och detta program gör det möjligt för oss att planera våra åtgärder ur en ny synvinkel och arbeta till förmån för kulturen på ett mer globalt , men också mer komplett och mer fördjupat sätt .
Jag gläds med er åt dessa tillfredsställande resultat som måste göra det möjligt för oss att , trots en budgetsituation som inte ligger i nivå med våra ambitioner , se framtiden an på ett mycket positivt sätt , och jag skulle vilja ta upp det som ordförande Gargani sade : kommissionen har gjort ett uttalande beträffande utvärderingen efter halva tiden .
Den har förklarat att i samband med den rapport den måste utarbeta i enlighet med artikel 7 i beslutet från parlamentet och rådet kommer den att genomföra utvärderingen av programmets resultat , och denna utvärdering kommer även att gälla de ekonomiska resurserna inom ramen för gemenskapens budgetplan .
Vid behov kommer rapporten att innehålla ett förslag till ändring av beslutet och allt detta före den 30 juni 2002 .
Mina damer och herrar , kära parlamentsledamöter !
Det är ett formellt åtagande , inte bara en mening på ett papper .
Allt detta måste leda oss till att stärka våra åtgärder till förmån för att lyfta fram ett gemensamt kulturområde , inom vilket våra kulturer kan utvecklas ytterligare i alla sina specifika karaktärer , all sin mångfald , men de kan också berikas ömsesidigt och övriga europeiska medborgare kan delta fullt ut .
Det är också tack vare parlamentet som vill att fler små åtgärder skall genomföras nära medborgarnas rötter snarare än stora spektakulära åtgärder .
Detta kommer att leda till att vi gör programmet " Kultur 2000 " till ett program för medborgarna .
Detta ökade deltagande från medborgarnas sida , som jag verkligen hoppas på , vill jag skall vara så brett och fruktbart som möjligt och jag förbinder mig att verka för att det blir en nåbar verklighet under de fem år som omfattas av programmet .
Jag vet att ni parlamentariker , i era regioner , i era länder , kommer att verka tillsammans med deltagarna i programmen för att alla dessa små blommor , som en kollega sade , skall bli en stor mångfärgad matta .
Jag skulle vilja att detta program blir en nåbar verklighet och att kulturen för våra medborgare utgör inte bara en berikande faktor , såväl på det personliga som det sociala och ekonomiska planet , utan även en rättighet som det handlar om att bekräfta , liksom ett tecken på en återfunnen sällskaplighet inom unionen .
Det är vad vårt europeiska program " Kultur 2000 " tillför .
Det är inte någon konkurrent till den kulturpolitik som bedrivs i de olika medlemsstaterna .
Den är nödvändig och jag skulle vilja se den utvecklas ytterligare .
Det är helt enkelt ett tillägg , ett komplement , ett byggande av en bro mellan de olika kulturerna i våra olika länder .
Att utvidga och berika de europeiska medborgarnas deltagande i kulturen förefaller mig alltså vara en grundläggande uppgift som motiverar våra ansträngningar och hur vi bör bedöma framgången med vår åtgärd och med vår union .
Flera parlamentariker har med rätta tagit upp det : om en union enbart består av ekonomi är den dödfödd .
Men om den består av kultur , om den består av civilisation , om den består av deltagande kommer den att bli levande .
Det är denna grund , mina damer och herrar , som jag har för avsikt att utveckla och jag kommer särskilt att ta hänsyn till följande inriktningar : för det första erbjuda möjligheter av innovativ karaktär för våra kreatörer så att deras talanger får det stöd de förtjänar i vårt program .
För det andra uppmuntra utbyte , rörlighet , utbildning inom kultursektorn .
För det tredje främja samarbete mellan kulturarbetare .
För det fjärde utöka allmänheten genom att bl.a. göra större plats för ungdomarna , och för det femte bevara och göra det gemensamma kulturarvet av europeisk betydelse mer känt , liksom de europeiska folkens historia .
Det nya programmet blir , genom sin struktur , sin organisation grundad på öppenhet , effektivitet och balans , det är jag säker på , ett instrument med lika hög prestanda som det blir grundläggande för våra åtgärder .
Fru talman !
Jag upprepar mitt tack till parlamentet för dess stöd och för att ännu en gång ha visat på den betydelse det fäster vid kulturen i unionssammanhang .
Jag är övertygad om att parlamentet inte kommer att bli besviket för att ha beviljat oss sitt stöd och jag förbinder mig att personligen successivt informera parlamentet om olika etapper i genomförandet av våra åtgärder , våra medborgares åtgärder , som jag hoppas skall bli stora åtgärder för unionens framtid .
Tack , fru kommissionär .
Jag tror att vi kan tacka vår föredragande ännu en gång .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.00 .
( Sammanträdet avslutades kl .
21.55 )
