 
Uttjänta fordon Nästa punkt på föredragningslistan är andrabehandlingsrekommendation ( A5-0006 / 00 ) från utskottet för miljö , folkhälsa och konsumentfrågor om rådets gemensamma ståndpunkt ( 8095 / 1 / 1999 - C5-0180 / 1999 - 1997 / 0194 ( COD ) ) inför antagandet av Europaparlamentets och rådets direktiv om uttjänta fordon ( föredragande Karl Heinz Florenz ) .
Herr talman , ärade damer och herrar , kära kolleger !
Årligen skrotas nio miljoner bilar i Europa .
Trots det faktum att dessa nio miljoner bilar inte längre kan köras har de den egenskapen att man handlar med dessa även mindre legalt även över gränserna , inte bara över gemenskapens inre gränser utan även över gränser som ligger utanför unionen .
Därför är det principiellt riktigt att Europeiska unionen upprättar allmänna spelregler för hur dessa nio miljoner fordon per år skall återvinnas och tas om hand .
Direktivet har enligt oss ett par svagheter som vi gärna vill rätta till här i kammaren genom ett direktiv som då verkligen blir framtidsinriktat .
Därför finns det en mängd ändringsförslag .
Jag personligen anser att man genom direktivets tillämpningsområde skjuter över målet .
Jag anser det inte nödvändigt att veteranbilar skall utgöra en del av direktivet .
Jag tycker heller inte att motorcyklar bör omfattas av direktivet , eftersom återanvändningen i fråga om motorcyklar är en så särskild kulturform att det inte behövs några europeiska direktiv för detta .
Inte heller för specialfordon eftersträvar jag nödvändigtvis höga återanvändningsnivåer .
Min önskan är den att specialfordon såsom ambulanser skall nå höga räddningsnivåer .
Det är mitt huvudsakliga bekymmer på det området .
Återvinningskraven på hur avfall från bilar skall hanteras i Europa föreskrivs efter mitt förmenande på ett bra sätt i direktivet .
Här kan det få stanna vid det som kommissionen har föreslagit .
Medlemsstaterna sörjer för att det finns motsvarande insamlingsanläggning där man tappar ur bilarna , tar hand om exempelvis över 32 miljoner spillolja , tömmer dem på bromsvätska etc .
En viktig komponent i direktivet är frågan : Vad vi skall göra med de gamla bildelarna ?
Vad gör vi med de skrotade produkterna ?
Man får inte blunda för att det kvantifierade målet är en viktig punkt när det gäller recycling ( återvinning ) och återanvändning ( recovering ) och vad det nu är , men det är inte den enda punkten .
För vi skall inte glömma : under en bils livscykel faller 80 procent av miljöbelastningen på körningen , 1 procent på sluthanteringen och 19 procent på tillverkningen av bilen .
Kvantifierade målsättningar är sålunda inte den enda parametern vid frågan om miljökonsekvenserna , utan en av många .
Jag är naturligtvis av den uppfattningen att vi behöver rigorösa mål .
Men kvoterna får inte bli ett självändamål , utan vi måste inse att helhetssynen på hur bilen belastar miljön är viktig .
Jag ser mycket hellre att vi kommer bort från en bil som i dag väger 1 400 kilo , som körs i genomsnitt i 200 000 km , till en bil som i framtiden väger endast 1 000 kilo och också körs i 200 000 km .
Trots allt skulle det då transporteras 400 kilo gånger 200 000 km mindre .
Detta är det sanna miljöpolitiska framsteget , för det leder till en kraftig minskning av koldioxid och detta är , om jag har förstått Kyotoprotokollet rätt , den viktiga beståndsdelen .
Därför tror vi att fordon som i framtiden på ett imponerande och påvisbart sätt använder sig av lättviktsmetoder producerar mindre koldioxid och ges speciella preferenser i förbränningskvoten .
Detta skall inte den enskilda medlemsstaten besluta om , utan det är ni , fru kommissionär , som tillsammans med er stab skall besluta om huruvida dessa lättviktsfordon - många talar även om 3-liter-bilar - skall erhålla speciella preferenser .
Vi är av den uppfattningen att det är riktigt .
Låt mig säga något om kostnaderna .
Vissa säger att tillverkarna borde få bära hela kostnaden - det skulle vara riktigt och mycket konsumentvänligt .
Detta kan man ifrågasätta mycket starkt , för tillverkarna kommer att lägga över alla kostnader på konsumenterna och tillägna sig ett återvinningsmonopol som borde vara statligt .
Jag kan bara varna er för att rösta för detta .
Det finns ändringsförslag som går ut på att kostnaderna skall delas , hälften åt tillverkarna och den andra hälften åt nybilsköparna .
Ur en sådan pool , ett sådant system , hur ni nu än föreställer er detta , kan man då från och med 2006 återta alla fordon i bilparken utan kostnad för den sista ägaren .
Detta är också min grupps uttryckliga önskan .
Vårt förslag om delning av kostnaderna har en alldeles avgörande fördel , nämligen att vi slipper bli domstolskandidat så snart vi har antagit direktivet .
För den återverkan som bilindustrin så listigt betalar tillbaka med är ett allvarligt problem som vi rimligen måste ta hänsyn till .
Därför föreslår jag att kostnaderna delas av den första ägaren och tillverkaren .
Förbud mot vissa material - naturligtvis behöver vi förbud mot vissa material .
Det finns farliga komponenter i bilen , dessa måste på sikt förbjudas .
Till det behöver vi ett instrument för påtryckningar .
Kommissionen har lagt fram några förslag som var för stränga , och vi har tagit fram alternativ till dessa .
Det finns en mängd bra ändringsförslag .
Parlamentet har fått större befogenheter .
Så låt oss utnyttja dessa !
Låt oss vara modiga nog att lägga fram och utveckla ett direktiv som pekar in i framtiden .
Ett direktiv som utvecklas endast för direktivens egen skull vore inte värdigt kammaren .
Jag ber om ert stöd .
Herr talman !
Jag får nästan lust att säga " puh ! " - äntligen har vi nått fram till andra behandlingen av det här direktivet , som har gett oss så mycket arbete , och givetvis enormt mycket för föredraganden , Florenz.Direktivet är enligt min mening inte alls tillfredsställande , eftersom det inte besvarar den verkliga frågan , nämligen vad man skall göra med redan övergivna fordon som i dag endast kan fraktas bort på samhällets och därmed skattebetalarnas bekostnad .
Man tillämpar således inte principen om att den som förorenar skall betala .
Redan övergivna fordon lämnas också i sticket av gemenskapens lagstiftning , eftersom de varken beaktas i texterna om avfallshantering eller i denna text om uttjänta fordon .
Direktivets enda förtjänst är att i det blickar man framåt .
Trots det har man inte löst problemet med de äldre bilar som används i dag , och som kostar mycket mer att återvinna .
Vi kan däremot ha en ganska stor tillförsikt inför framtiden med tanke på vilka insatser biltillverkarna är beredda att göra , å ena sidan för att finna material som är lättare att återvinna och å andra sidan för att få igång återvinningsprocessen .
Jag vill också insistera på det faktum att vi måste behålla en flexibilitet mellan återvinning , återanvändning och förbränning när det gäller de nya särskilt lätta material som kan dämpa bilkonsumtionen , och därmed utsläppen .
Detta är ett problem som handlar om förenligheten mellan våra direktiv om uttjänta fordon och de äldre direktiven , bl.a. fordons- och oljeprogrammet , som vi röstade igenom för några år sedan .
Man kan således glädjas åt att utskottet för miljö , folkhälsa och konsumentpolitik har varit förnuftigt och infört ett undantag för de veteranbilar som utgör en del av vårt industri- och kulturarv - så att det inte skall råda något tvivel om den saken .
Sammanfattningsvis är direktivet inte tillräckligt ambitiöst för att problemen med den nuvarande bilparken skall kunna lösas .
Det är dessutom ganska så hycklande vad gäller de vrak som fortfarande belamrar våra skogar , sjöar och parker .
Återigen , principen att den som förorenar skall betala tillämpas inte , och det är alltid skattebetalarna som får stå för notan .
Herr talman , fru kommissionär , kära kolleger !
När man ser de flygblad som har delats ut under de senaste veckorna så tror man att det är en möjlig miljökatastrof eller den europeiska bilindustrins död vi diskuterar här. inte något av detta stämmer .
Vi måste se med nyktra ögon på att direktivet som ligger framför oss på bordet är ett bra direktiv .
Det innebär miljömässiga framsteg för Europa , och vi kan vara stolta om vi kan få till stånd och förankra direktivet i lag .
Förvisso , det finns en punkt som vi är oense om .
Med tanke på direktivets dimensioner är det måhända en liten punkt , men det är detta oenigheterna handlar om .
Det gäller frågan om kostnaderna för återvinningen .
Här skiljer vi oss i väsentliga delar från diskussionen i rådet förra året .
Där drogs nämligen kostnadsbefrielsen för sista ägaren och frågan om finansieringen över en kam , och kostnadsbefrielsen för sista ägaren ifrågasattes .
Vi här i kammaren fattade entydigt beslut i februari förra året - och detta stöder vi , just vi socialdemokrater - kostnadsbefrielsen för sista ägaren är för oss odiskutabel !
Men vem betalar för de fordon som skall skrotas och tas om hand ?
För oss är det självklart att tillverkaren skall göra detta vad gäller nya bilar , därför att detta också är ett incitament för tillverkaren att ta fram och tillverka återvinningsvänliga bilar .
Men vad händer med fordonen som rullar på gatorna ?
Ett exempel : Firman Rover i Storbritannien skulle , om man blev ansvarig för alla uttjänta fordon , bli ansvarig för 5,8 miljoner bilar i Europeiska unionen och omgående tvingas öronmärka 250 miljoner euro för att spara ihop till återvinningskostnaderna , medan en tillverkare av liknande bilar från Korea behöver lägga undan ett peanuts-belopp - som en företrädare för Deutsche Bank en gång uttryckte det .
Här finns en snedvridning av konkurrensen som inte har med miljöskyddet att göra utan enbart inverkar på investeringsförmågan , och på arbeten för de människor som bygger bilar här i Europa .
I så måtto föreslår jag att en fond för de gamla fordonen bildas , ur vilken återvinningskostnaderna för de uttjänta fordonen sedan betalas så att principen om kostnadsbefrielse säkras .
Jag kan förstå att kolleger från länder utan biltillverkning säger ja , tillverkarna skall betala alltihop , och problemet med snedvridningen av konkurrensen genom öronmärkta reserver intresserar oss inte !
Men jag ber dessa kolleger visa solidaritet med de drygt två miljoner människor som tillverkar bilar i Europa , som på så sätt finansierar sina liv , så att dessa arbetsplatser kan garanteras även i framtiden .
Jag är för stränga miljökrav , det vet ni från Auto / Oil-programmet och diskussionen om gränsvärdena för avgaser .
Men jag anser att kraven måste vara lika för alla !
Herr talman , herr kommissionär , kolleger !
Jag tror att vi behöver detta direktiv .
För det första eftersom det innehåller en tydlig beskrivning av miljömålsättningarna .
För det andra eftersom detta direktiv kan stimulera återanvändning , och det är viktigt .
För det tredje finns det ett tydligt tillvägagångssätt för att motverka föroreningen från tunga metaller .
Det är också en viktig punkt .
Direktivet ger en europeisk ram , bland annat också för medlemsstater som redan har ett system och som vill fortsätta att arbeta med det systemet .
Vi måste således i första hand bibehålla procentandelarna i fråga om återvinning , för därigenom uppmuntrar man naturligtvis teknisk förnyelse och olika sätt att hitta en lösning för material som vi ännu inte riktigt vet vad vi skall göra med .
För det andra måste vi låta de omständigheter som står i den gemensamma ståndpunkten vara oförändrade .
Så från och med år 2006 gäller kostnadsfri inlämning för alla bilar , kostnadsfri för den sista ägaren .
Det är naturligtvis helt klart en mycket viktig punkt .
Den får vi inte tumma på .
Är detta en för stor börda ?
Det finns dock en sak som vi inte får glömma bort .
Direktivet handlar om fullständiga bilar , alltså bilar där inga viktiga delar saknas .
Enligt experterna är det inte många av dessa fullständiga bilar som är värdelösa .
För återvinning , återanvändning av delar , det är en sektor som inte nödvändigtvis är förlustbringande .
Tvärtom , det finns för närvarande ett stort antal företag som lever av detta och som därigenom utan problem kan förtjäna sitt levebröd .
Detta direktiv stimulerar hela denna sektor .
Det handlar om en sektor som utgörs av små och medelstora företag .
Eftersom transportkostnaderna i detta fall ligger på en hög nivå måste det också bli fråga om ett starkt decentraliserat system , för att flytta ett vrak mer än 100 kilometer är inte någon lönsam verksamhet .
Jag tycker att det är en bra idé att detta direktiv inte skall gälla för historiska bilar , och jag anser att det måste vi lägga till .
Så enligt min uppfattning bör veteranbilar befrias från detta .
Det är också bra att vi tydligt lägger ansvaret hos producenten .
Det är en grundläggande princip och den måste vi hålla fast vid .
Han är ansvarig för konstruktionen .
Han kan således göra en mycket stor insats för miljön i samband med denna konstruktion .
Vi måste också hålla fast vid att kostnaderna skall bäras av producenten , helt eller till övervägande delen , vilket står i den gemensamma ståndpunkten .
Jag anser att det är en balanserad princip som inte utesluter några andra saker .
Min uppfattning är att vi måste behålla denna .
Därför kommer vår grupp att stå kvar så nära den ursprungliga gemensamma ståndpunkten som möjligt och inte förändra denna ståndpunkt på de väsentliga punkterna .
För vi vet naturligtvis allesammans att det var mycket mödosamt att få till stånd denna ståndpunkt i rådet , att det var en svår balansövning att uppnå denna gemensamma ståndpunkt .
Vi får , enligt min uppfattning , från vår sida inte sätta denna gemensamma ståndpunkt i fara , för detta är ett direktiv som vi absolut behöver av miljöskäl .
Jag uppmanar er att stödja denna gemensamma ståndpunkt .
Vår grupp kommer i vilket fall att göra detta i så stor utsträckning som möjligt av miljöskäl eftersom vi har detta direktiv och eftersom det är ett balanserat direktiv som innehåller en mängd saker , en mängd invändningar , till exempel i fråga om kostnadsfördelningen .
Herr talman , kolleger !
I dag har vi ett viktigt beslut att fatta .
Stöder Europaparlamentet den ekologiska principen om producentansvar , det vill säga att fordonstillverkarna har ansvaret för bilar när de har blivit bilvrak ?
Nej , säger kristdemokraterna i ändringsförslag 38 : fordonstillverkare och bilister skall dela kostnaderna lika .
I förpackningsdirektivet , där denna kompromiss om att dela lika står , kan man se att detta inte fungerar .
Förpackningar är fortfarande ett stort nedskräpningsproblem i Europa och en belastning på miljön .
En del av socialisterna under ledning av Bernd Lange säger : " Ja , den här principen är bra , men vi skall inte införa den förrän år 2010 eller år 2012 enligt ändringsförslag 45 . "
I den gemensamma ståndpunkten står det år 2006 .
Enligt Gruppen De gröna ger det bilindustrin mer än tillräckligt med tid att förbereda sig .
Jag uppmanar därför mina kolleger att inte stödja kristdemokraternas ändringsförslag 38 och 45 av ett antal socialister .
Om fordonstillverkarna själva måste stå för kostnaderna för återvinning av sina bilar , då kommer de att konstruera dem så att de blir lättare och billigare att återanvända .
Då kommer problemet med plast , PVC , att försvinna från bilar och ersättas av bioplast framställd av växter .
När allt kommer omkring är det billigare , också för konsumenterna .
I tjugo års tid har en majoritet i parlamentet försökt att göra den europeiska miljöpolitiken grönare .
I dag hotar denna gröna position att gå förlorad under tryck från framför allt den tyska och franska bilindustrin .
Därför , kolleger , rösta emot ändringsförslagen 38 och 45 .
Vi i Gruppen De gröna stöder i stora drag den gemensamma ståndpunkten .
Herr talman !
Avfallet från uttjänta bilar är ett av våra riktigt stora miljöproblem , både vad gäller avfallsmängd och utsläpp av miljöskadliga ämnen .
Vi i GUE / NGL-gruppen vill därför ha ett så heltäckande och konsekvent regelverk på området som bara är möjligt .
Med detta direktiv har vi en möjlighet att ta ett stort steg framåt , men det förutsätter att rådets ståndpunkt inte trasas sönder och försvagas i parlamentets behandling .
Flera av de ändringsförslag som har lagts fram skulle , om de antogs , försvaga direktivet mycket kraftigt .
Det gäller framför allt ändringsförslag från PPE-gruppen , men tyvärr också några ändringsförslag från Lange , som jag ser det .
Det är inte svårt att ana att vissa länders bilindustri , t.ex. den tyska , har utfört ett ganska hårt lobbyarbete inför antagandet av detta direktiv .
För oss är det avgörande att följande principer skall gälla : Förorenaren skall betala .
Det innebär att det är tillverkaren som skall ta det fulla ansvaret också ekonomiskt för återvinning av fordonen .
Det måste finnas regler även för befintliga fordon .
Vad gäller det kan vi inte godta att rådets ståndpunkt vad gäller datum för ikraftträdande skulle försvagas .
Procentsatserna och kraven på återvinning vid vissa årtal får inte försämras .
Dessutom är det viktigt att begränsa användningen av farliga ämnen som bly .
Vi kommer att rösta emot alla ändringsförslag som går i motsatt riktning i förhållande till detta .
Om de ändringsförslag skulle antas som kraftigt försvagar direktivet , vore det mycket negativt , inte bara ur miljösynpunkt utan också för Europaparlamentets trovärdighet i miljöfrågor .
Det hänvisades tidigare i debatten till att man skall tänka på de miljoner människor som arbetar i bilindustrin i olika länder och de länder som har en stor bilindustri , t.ex. mitt eget hemland Sverige .
Jag har själv varit bilarbetare innan jag blev invald .
Jag tror mig vara en av få i detta parlament som har stått vid ett löpande band och monterat bilar .
Jag tycker att man skall ställa mycket hårda krav på bilindustrin .
Det gynnar nämligen de moderna biltillverkarna som tänker miljövänligt och går snabbt framåt .
Det är precis den typ av bilindustri som vi skall uppmuntra i Europeiska unionen .
Herr talman !
Det gläder mig mycket att parlamentet nu prioriterar miljöskyddet , vilket medborgarna i Europa med all säkerhet också gör .
Det råder inget tvivel om , att övergivna bilar utgör ett allvarligt hot mot den visuella och fysiska miljön .
Våra medborgare förväntar sig i detta hänseende att vi skall bevaka deras intressen .
Varje år skrotas mellan 8 och 9 miljoner fordon inom Europeiska unionen .
Detta genererar i sig en stor mängd avfall .
Biltillverkare , underleverantörer och tillverkare av utrustning måste anstränga sig för att begränsa användningen av farliga ämnen och måste därför i planeringsskedet se till att återanvänt material kan användas i tillverkningen av bilar .
Vi vet att det i Nederländerna finns auktoriserade behandlingscentraler som samlar upp uttjänta fordon , och denna metod bör spridas över hela Europeiska unionen .
Sett ur ett irländskt perspektiv vet jag att det irländska miljödepartementet redan har börjat samråda med företrädare för motorindustrin för att se till att lämpliga uppsamlingsplatser upprättas inom en snar framtid för att ta hand om uttjänta fordon på Irland .
Jag ser inget skäl till varför man inte skulle kunna organisera ett tillståndssystem för uppsamlingsplatser över hela Europa , för att skrota de 8 till 9 miljoner fordon som man årligen gör sig av med inom Europeiska unionen .
Biltillverkare skall lämna information om hur stor del av de begagnade bilarna som kommer att kunna återanvändas , återvinnas och återställas under de kommande åren .
I enlighet med de nya bestämmelserna i Amsterdamfördraget har samtliga 370 miljoner konsumenter inom Europeiska unionen rätt till konsumentrelaterad information .
Jag tror att EU : s konsumenter kommer att stödja de biltillverkare som tillämpar de miljövänligaste metoderna under det kommande året .
Den sista frågan jag vill ta upp är att man i bestämmelserna och lagstiftningen måste ta hänsyn till den traditionella bilsektorns speciella ställning i hela den Europeiska gemenskapen , på grund av den roll denna har i förhållande till den sociala sektorn samt mot bakgrund av miljömässiga och ekonomiska hänsynstaganden .
Herr talman , ärade ledamöter !
Direktivet om uttjänta fordon är verkligen en milstolpe på vägen mot en bättre miljö i detta vårt Europa .
Det verkar också som om man verkligen har ansträngt sig för att komma fram till en intelligent återanvändning av materialen , en minskning av det förorenande avfallet och ett främjande av tekniska innovationer .
Vad detta beträffar är vi verkligen på rätt väg men , som några kolleger redan har betonat , är det reella problemet möjligheten att tillverkarnas ansvar blir ett solidariskt ansvar .
Jag skulle vilja säga att man i Italien har tagit betydande steg framåt på detta område .
Vi var kanske först i Europa med att införa ett regelverk som uppmuntrar till att ta uttjänta fordon ur bruk , men vi har också i vårt land en ganska gammal bilpark och därmed allvarliga bekymmer för de marknadsproblem detta direktiv skulle kunna medföra .
Jag tror att man måste analysera fenomenet på allvar .
I Italien har man kommit till en inlämnings- och återvinningsgrad på omkring 80 procent , men det finns ett marknadsproblem som skulle kunna orsaka en smärre kris vad sysselsättningen beträffar .
Eftersom vi i Italien har en industri som ofta tillgriper tillfälliga och permanenta friställningar kan detta medföra allvarliga svårigheter för löntagarna i olika delar av landet .
Jag märker att parlamentet ibland är litet extremistiskt och intar ståndpunkter som antingen är ytterligt gröna eller raka motsatsen .
Därför tycker jag att man borde försöka förena de två kraven och finna en syntes .
Florenz och andra ledamöter verkar ha funnit den och försöker när allt kommer omkring förena de två åsikterna .
Resultatet är dessa intressanta ändringsförslag .
Här tror jag att man kan hitta en avvägd lösning på problemet , det vill säga att förena miljökraven med marknadens och sysselsättningens behov .
Herr talman !
Detta direktiv behandlar det förhållandevis lilla men växande problemet med övergivna bilar samt frågan om en mera strukturerad skrotning av uttjänta bilar .
I den utsträckningen kan det tänkas vara önskvärt , trots att det inte är något brådskande ärende .
Huvudfrågorna är nu vem som betalar 262 euro per bil för de 9 miljoner bilar som skrotas varje år .
Vem betalar för uppsamlingen , demonteringen , skrotningen och så vidare ?
Och skall direktivet retroaktivt omfatta varje bil som någonsin tillverkats ?
Kommissionens förslag , den allmänna ståndpunkten , är att tillverkarna skall betala allt .
Detta skulle betyda miljarder pund eller euro för vart och ett av de större företagen i varje land inom Europeiska unionen .
Denna kostnad skulle ofrånkomligen föras över på priset och följaktligen på de nya bilarnas köpare .
Eftersom europeiska biltillverkare har verkat här under många fler decennier än företag från Japan , Korea och andra länder , skulle det ligga till mycket större last för de äldre europeiska företagen och utgöra en konkurrensfördel för deras konkurrenter från andra länder .
Jag uppskattar Florenz , Lange och andra som från partisplittringens båda sidor försökt uppnå en kompromiss baserad på delade kostnader .
Jag rekommenderar också det ändringsförslag som jag undertecknat samt uppmanar mina kolleger från Tyskland , Italien , Irland , Spanien , Sverige och Storbritannien att eliminera denna åtgärds retroaktiva drag .
Retroaktiv lag är dålig lag , den är ofta orättvis och ofta ogenomförbar .
De flesta demokratiska parlament i den fria världen förkastar den av princip såvida det inte föreligger ett överväldigande offentligt intresse , vilket det tydligen inte gör i det här fallet .
Det är därför jag har manat till en omröstning med namnupprop om detta .
Vi kan då se vem som är beredd att rösta för retroaktivitet med tvivelaktig legalitet , vilket skulle innebära en kostsam belastning för varje framtida bilköpare och ett förödande slag mot den europeiska bilindustrin .
Herr talman , mina kära kolleger !
Jag vill än en gång helt kort påminna om vilka ekonomiska frågor som står på spel med detta direktiv , och förnya mitt stöd till de ändringsförslag som min kollega Bernd Lange har ingivit .
Fördelen med dessa ändringsförslag - jag vill insistera på detta - är att de sammanjämkar miljökrav och ekonomiska absoluta krav .
Rådets gemensamma ståndpunkt innebär att biltillverkarna skall stå för hela eller en avsevärd del av kostnaderna för återtagande och återvinning av fordon .
Men som Lange så väl uttryckte det : för de europeiska tillverkarna är den lösningen fullkomligt orättvis .
Eftersom jag kommer från ett land där det faktiskt finns biltillverkare , kan jag tala om att det är en omöjlighet att retroaktivt ålägga dem ett totalt finansiellt ansvar för alla de fordon som kommer från deras fabriker och som nu rullar på vägarna , vilket innebär ett ansvar för kostnader som ålagts 80 procent av den europeiska bilparken .
Denna lösning är oacceptabel , eftersom tillverkarna inte har kunnat integrera miljökraven i sina tillverkningsprocesser och självkostnadspriser , de miljökrav som vi ålägger dem i dag .
Den gemensamma ståndpunkten sätter de europeiska tillverkarna i ett ofördelaktigt läge gentemot de tillverkare som nyligen trätt in på den europeiska marknaden .
Vi är självklart inte här för att försvara det ena eller andra nationella intresset eller den ena eller andra industrilobbyisten .
Vi är däremot här för att bygga upp ett Europa som kan konkurrera på världsmarknaden och för att försvara sysselsättningen inom de ekonomiska sektorer där vi faktiskt är konkurrenskraftiga .
Av det skälet , kära kolleger , ber jag er att stödja de ändringsförslag som ingivits av Bernd Lange och som kommer att stödjas av Europeiska socialdemokratiska partiets grupp .
Faktum är att dessa ändringsförslag förlikar samtliga intressen - ekonomiska intressen och miljökrav - samtidigt som medlemsstaterna förblir fria att besluta om de närmare bestämmelserna för genomförandet av dessa krav , eftersom de system som nu gäller i medlemsstaterna - och det finns de som fungerar helt tillfredsställande - enligt förslagen skall få finnas kvar i fortsättningen .
Herr talman , fru kommissionär !
Det förslag till direktiv om uttjänta fordon som vi i dag ägnar oss åt syftar dels till att garantera ett starkt miljöskydd inom unionen , och dels till att säkra en fortsatt väl fungerande inre marknad för denna sektor .
Jag vill bara kort säga att historiska bilar och veteranbilar givetvis skall undantas från tillämpningsområdet för detta direktiv .
Vi är väl alla överens om att bilarna också utgör en del av vårt kulturarv .
En av stötestenarna avser artikel 12 , dvs. när direktivet skall börja tillämpas .
Parlamentets föreslagna lösning , nämligen 18 månader efter det att direktivet trätt i kraft för nya bilar , är föga realistiskt .
Den europeiska bilparken omfattar tiotals miljoner bilar som skall återtas utan att de har tillverkats för att återvinnas .
Den gemensamma ståndpunkten var mer praktisk , eftersom den fastställde år 2006 för de bilar som redan är i trafik .
Detta skulle dessutom ge företagen tid att uppbringa resurser för att hantera de tillkommande kostnaderna .
I likhet med min grupp kommer jag således att stödja den gemensamma ståndpunkten , som förefaller vara en balanserad kompromiss mellan företagens begränsningar och nödvändiga framsteg på miljöskyddsområdet .
Herr talman , kära kolleger !
Europaparlamentet står i dag inför ett viktigt beslut .
Skall vi arbeta för ett framtidsorienterat miljö- och konsumentskydd eller skall parlamentet , vilket man kan befara enligt ändringsförslagen från Florenz , Lange och andra , göra sig till bödelsdräng åt den tyska bilindustrin ?
Parlamentets trovärdighet som en av pionjärerna för miljöskydd står på spel .
Det vore mer än genant om Europaparlamentet skulle urvattna det som regeringarna i de 14 medlemsstaterna och Europeiska kommissionen har beslutat vad gäller tillverkaransvaret och skyddet av miljön !
Den avsikt Florenz och Lange har med ändringsförslagen är tydlig : direktivet skall förstöras !
Genom det föreslagna delade ansvaret skall principen om att förorenaren skall betala urholkas och produktinnovationer undergrävas .
Genom uppbyggnaden av talrika hinder vill de ingenting annat än att förhindra en effektiv ekologisk politik för avfallsströmmar , och via typgodkännanden vill de fördröja tillämpningen av direktiven med tolv år eller mer .
Detta är fullkomligt oacceptabelt .
Jag vädjar därför alldeles särskilt till de tyska ledamöterna : Förhindra att det i dag uppstår en stor politisk skada !
Den rödgröna förbundsregeringen har inte precis skördat några större lagrar i debatten om direktivet för uttjänta fordon .
Låt inte detta fortsätta !
Det ständiga gnället om konkurrensnackdelen är löjeväckande när det egentligen bara handlar om en konkurrensnackdel för den tyska bilindustrin .
Var företrädare för folket , och låt er inte degraderas till företrädare för Volkswagen !
Rösta för miljö- och konsumentskyddet och för innovationer i bil- och återvinningsindustrin !
Herr talman !
Vi har diskuterat detta direktiv sedan 1997 .
Nu är det dags att vi kommer fram till en överenskommelse .
Eftersom jag mer eller mindre delar de åsikter som min kamrat Sjöstedt och De grönas företrädare De Roo framförde , tänker jag inte använda de två minuter jag har till mitt förfogande utan bara betona två frågor .
För det första , och det är kanske det viktiga i förslaget : tanken både angående återvinning och återanvändning om att man skall använda material som är mindre förorenande .
En annan viktig punkt är att avfall inte skall brännas eller sönderdelas , men inte bara när det gäller det som innehåller bly , kadmium och kvicksilver utan också det som innehåller PVC .
Vi diskuterar denna fråga i ett annat forum i parlamentet .
Den andra frågan gäller vem som skall stå för kostnaderna .
Jag håller med de tidigare talarna när de säger att den som förorenar skall betala , och det har aldrig sagts bättre tidigare än i detta förslag .
Tillverkarna skall betala , även om vi alla vet att kostnaderna i slutändan kanske läggs på konsumenterna , och de skall ta hand om kostnaderna före 2006 så som föreslås i vissa ändringsförslag .
Vi instämmer mer med ändringsförslaget från första behandlingen .
Det är också viktigt att fastställa en viss procent och det datum då fordonen skall bestå av återvinningsbart material .
Jag tycker att man enligt förslaget förlitar sig på alltför långa tidsfrister .
Slutligen , herr talman , anser jag att det är nödvändigt att gynna små och medelstora företag som , efter sträng kontroll och erhållande av vederbörliga tillstånd , kan skapa sysselsättning i detta så viktiga arbete , och på så sätt undvika storföretagens monopol .
Herr talman , kära kolleger !
I dag måste Europaparlamentet åta sig ett verkligt ansvar .
Det handlar om vad vi skall göra med de miljoner fordon som vi överger varje år .
I vissa av våra stater har frivilliga miljöavtal redan tecknats för att våra diken , kanaler och fält inte längre skall fyllas av anskrämliga och farliga vrak , som en och annan skrämd höna har flytt .
Jag kommer från ett land som är stolt över sin bilindustri och dess kommersiella framgångar , såväl i Europa som i tredje land .
Mitt lands internationella nimbus är en mätare på dess betydelse .
Jag känner till den europeiska bilindustrins aktiva beteende ; den har satt igång ett omfattande forskningsprogram i syfte att upprätta ett nationellt informationssystem för nedmontering av gamla fordon .
Jag är medveten om vilka svårigheter rådet har stött på för att finna en kompromiss .
Därför måste vi i dag vara alkemister med förståelse och omsorg om vår miljö .
Detta sekel kommer att bli avfallshanteringens sekel , i annat fall blir det inget sekel alls .
För min del bör man tillämpa principen att den som förorenar skall betala .
Jag är säker på att bilindustrin , som visar en ständigt större respekt för miljön , har förväntat sig en sådan insikt .
Den tar dessutom sitt ansvar .
Men det åligger staterna att genomföra detta direktiv , och vi får akta oss för att göra det alltför detaljerat , eftersom de industriella traditionerna , nedmonterings- och skrotningsprocesserna ser olika ut beroende på om man är i Italien eller Finland .
Jag motsätter mig det faktum att bilägarna skall göras ansvariga .
Alla dessa kvinnor och män som rör på sig överallt i Europa , de betalar sin bil , sin nationella skatt , sin katalysator , sin bränsleskatt - de betalar således redan ett mycket högt pris för denna fantastiska maskin och friheten att förflytta sig .
Det skulle vara väl oförsiktigt - av mina kolleger i de stora grupperna med federalistisk böjelse - att vilja göra Europaparlamentet så impopulärt genom att kunna tänka sig ett delat ansvar mellan ägaren och tillverkaren .
Hur skall man dessutom kunna skapa en fond för att betala fordonsåtervinningen och förvaltningen av inomeuropeiska operationer ?
Vem kommer att betala återvinningen av min bil som jag köpt i Frankrike om jag låter registrera den i Belgien ?
Vilken nationell fond kommer att ta på sig ansvaret för mitt uttjänta fordon ?
Vi får också akta oss för att oroa företagarvärlden med den rättsliga osäkerhet som har att göra med en oacceptabel retroaktivitet .
Det är inte vår sak , här , att i dag dra igång en vedergällningsaktion med stöd av lagstiftning , vi bör i stället fortsätta på vår väg genom att förorda en hållbar utveckling .
Herr talman !
Europaparlamentet med utskottet för miljö , folkhälsa och konsumentfrågor i täten föresätter sig mestadels att kritiskt bedöma förslag från Europeiska kommissionen eller rådet och förbättra dem från miljösynpunkt .
Nu hotar en gedigen gemensam ståndpunkt från rådet att här i parlamentet bli sämre från miljösynpunkt .
Varje år skrotar vi ett stort antal bilar med många farliga ämnen .
Därför är förebyggande åtgärder med avseende på avfallsämnen viktiga .
Vi bör också sträva efter så små mängder som möjligt av tungmetaller och andra farliga ämnen och material .
Dessutom bör biltillverkarna ta hänsyn till att dessa bilar tillverkas på ett sådant sätt att det är enkelt att demontera och återanvända dem .
Resterna av bilvraket kräver också en adekvat behandling .
Jag stöder därför helhjärtat de procentsiffror för återanvändning och återvinning som föreslagits av rådet .
Numera är det ekonomiskt möjligt att genomföra en fullständig demontering av bilvrak .
Detta innebär att vi överger sönderdelning av bilvrak .
De uppställda målen är säkert genomförbara , och i Nederländerna har återvinningen redan uppnått ett värde på 86 procent .
Det bästa sättet att sörja för en god insamling är att den sista användaren kan lämna in bilen utan kostnad till en auktoriserad behandlingsanläggning .
Kostnaderna för behandlingen kan sedan tas ut på priset för nya bilar .
De förslag som lagts fram av vissa parlamentsledamöter skadar detta system på ett allvarligt sätt .
Det så kallade delade ansvaret är mycket opraktiskt och stimulerar inte till någon innovation .
Om systemet med kostnadsfri inlämning tillämpas kommer det också att visa sig att kostnaderna för behandling kommer att sjunka avsevärt .
Slutligen måste detta direktiv träda i kraft så snabbt som möjligt .
Ett segdraget förlikningsförfarande innebär en onödig försening som går ut över miljön .
Låt oss vara nöjda med den gemensamma ståndpunkt som nu föreligger ; då behöver vi inte göra någonting annat än att komplimentera och lyckönska rådet till det uppnådda resultatet .
Herr talman !
Jag vill ge kollega Florenz ett stort erkännande .
Han har under tryck , inte bara från sina kolleger utan också från bilindustrin , gjort ett gott arbete .
Lägg därtill att Florenz också var tvungen att göra detta med sin ekologiskt gröna inställning , var tvungen att mot den bakgrunden finna en kompromiss , och det var inte lätt .
Allmänt sett är jag inte missnöjd med den gemensamma ståndpunkt som här ligger framför oss , och i vilket fall som helst inte med den filosofi som ligger bakom den gemensamma ståndpunkten .
Det är två punkter som jag skulle vilja säga något om .
Det gäller veteranbilarna och motorcyklarna , vilka mycket riktigt skall undantas från direktivet , och den andra punkten är hela den kontroversiella frågan om vem som egentligen bär ansvaret för återtagandet av bilarna .
Jag vill inte tumma på texten i den gemensamma ståndpunkten .
Producenten är ansvarig , måste vara ansvarig , och slutanvändaren måste utan kostnader kunna återlämna bilen .
Jag tror att det finns för mycket ogrundad rädsla .
Billobbyn har fört för många bakom ljuset .
Jag vill därför än en gång säga till kollegerna att erfarenheterna visar att kostnaderna för denna behandling läggs på priserna .
Det är inte så höga kostnader .
I den medlemsstat som jag kommer ifrån handlar det om 150 gulden per bil .
Det innebär att man börjar på dag noll , och man kan då också behandla de gamla bilarna direkt .
Då kan också en mycket stor industri direkt byggas upp som innebär att man ser till att de bilkyrkogårdar som tidigare var en vanlig syn i våra medlemsstater upphör att existera .
Jag vill alltså inte tumma på den punkten i kompromissen .
Jag tror att det är bra att vi så snabbt som möjligt sinsemellan godkänner den lagstiftning som nu ligger framför oss .
Det är bra , eftersom det innebär att de nio miljoner bilar som varje år kommer ut på vägarna i Europa också tas om hand på ett ordentligt sätt .
Det kommer oss allesammans till godo .
Herr talman !
Det föreliggande direktivet är en viktig åtgärd för att förebygga att vi får farligt avfall från uttjänta fordon , och det är viktigt för att främja återanvändning och återvinning av material från skrotade bilar .
Jag menar därför att det är miljömässigt avgörande att förbudet mot att använda giftiga tungmetaller genomförs fullt ut , och att vi inte försvagar tillverkarnas ansvar .
Gör vi detta tar vi bort incitamentet för tillverkarna att konstruera och tillverka bilar som ger mindre avfall .
Det gemensamma systemet som efter mycket bekymmer antogs av rådet , som kommissionen stöder , och som också stöds av parlamentets utskott för miljö , uppfyller fullständigt de fastställda miljökraven och jag tycker därför att det är mycket egendomligt och oförståeligt att se ändringsförslag från ledamöter av utskottet för miljö som syftar till att väsentligt minska biltillverkarnas ansvar .
Om dessa ändringsförslag antas , menar jag att parlamentets trovärdighet i miljöfrågor allvarligt måste ifrågasättas .
Vi i parlamentet har hittills varit en positiv katalysator för miljöskydd och nu blir vi en negativ miljöfaktor i denna fråga i Europa , om ändringsförslagen från Florenz och Lange antas .
Om vi dessutom försvagar tillverkarnas ansvar i denna fråga , kommer det att få allvarliga konsekvenser för senare frågor på andra områden , t.ex. det kommande direktivet om elektronik- och datorskrot .
Jag vill därför gärna uppmana parlamentets ledamöter att vi utan hänsyn till grupptillhörighet röstar emot alla de ändringsförslag till den gemensamma ståndpunkten som kommer att försvaga den miljömässiga standarden och som kommer att minska tillverkarnas ansvar .
På så sätt kan vi uppnå ett miljömässigt anständigt resultat .
Herr talman !
Detta förträffliga direktiv kommer att göra slut på dumpandet av gamla bilar , gynna återvinningen och framför allt uppmuntra tillverkarna att utforma bilar som lätt kan återvinnas .
Men vem skall stå för kostnaderna ?
Vilket system som än införs , kommer kostnaden slutligen att föras över på konsumenten .
Det bästa sättet för oss att uppnå våra miljömål är att göra tillverkarna till vårt verktyg såväl för insamlingen av pengarna som för skrotningen och återvinningen av bilarna .
Tillverkarna har lurat Florenz och Lange att lägga fram ändringsförslag här som allvarligt försvagar dessa förslag .
Låt er inte luras av biltillverkarna !
Om ni vill dra full nytta av detta direktiv , använd er röst till att förkasta dessa ändringsförslag .
Herr talman , fru kommissionär , kära kolleger !
I motsats till vad vi skulle kunna tro är denna debatt inte av teknisk art .
Den har blivit högst politisk .
I går hedrade vi vår institution med en politisk debatt - vi skulle vanhedra oss själva om 314 ledamöter i dag gav efter för vissa biltillverkares lobbygrupper .
Genom att begära att konsumenterna skall stå för hälften av kostnaderna för återtagande av uttjänta fordon , vilket ändringsförslag 38 föreskriver , samtidigt som den gemensamma ståndpunkten kräver att tillverkaren skall ansvara för hela återtagandet , skulle Europaparlamentet för första gången inte framträda som en garant för försvaret av de europeiska konsumenterna och medborgarna , utan i stället bli något av en resonanslåda för lobbygrupperna .
Det kan vi inte acceptera .
Det skulle vara ett prejudikat som öppnade dörren för alla slags påtryckningar inom många andra områden .
Det skulle också vara första gången som Europaparlamentet försvagade rådets ståndpunkt , när vi i allmänhet kritiserar rådets ståndpunkter för att inte räcka till .
Ett system för gratis återtagande av gamla fordon och ett utökat antal fordon som skall återvinnas är exempel på åtgärder som kommer att få såväl återvinningsverksamheten som den därmed förknippade sysselsättningen att växa .
Med tanke på konsumenterna , miljön och de nya arbetstillfällen som kan skapas inom återvinningssektorn , får vi absolut inte ändra rådets gemensamma ståndpunkt , som i sin nuvarande version är helt godtagbar .
Herr talman !
Liksom så många andra här i dag tror jag att detta är en bra åtgärd .
Det är en nyttig åtgärd och nödvändig för oss alla .
De flesta tekniska frågorna är lösta .
Det återstår att slutgiltigt godkänna vissa detaljer , men de flesta tekniska frågorna är lösta .
Vi har kommit fram till den sista frågan .
Under debatten vid den första behandlingen var det endast utskottet för ekonomi och valutafrågor som ställde den här frågan och det var bara jag själv i egenskap av den som författat utskottets yttrande som ställde den frågan i parlamentet .
Den är mycket enkel : Vem betalar ?
Kommissionens allmänna ståndpunkt innebär en rimlig kompromiss på så sätt att tillverkarna skall betala en betydande del av kostnaden , inte hela kostnaden som Bowis nämnde av misstag .
I själva verket så litet som 20 procent eller en femtedel av kostnaderna , enligt juristerna .
Detta är inte orimligt .
Om man ser på konsumenten i Storbritannien som köper en Rover , som Lange pekat på , eller vilket annat bilmärke i Storbritannien som helst för den delen och som i åratal har betalat överpriser för dessa bilar , långt över jämförbara priser i andra delar av Europa , varför skall de betala ?
De har redan betalat .
Varför skulle de här människorna , som skattebetalare eller som framtida bilköpare , åter betala för skrotning av ett fordon som tillverkaren har gjort vinst på ?
Jag kan inte acceptera det .
Enligt vissa ändringsförslag här i dag föreslås det att detta bör vara fallet .
Jag kan inte acceptera det och jag kommer inte att rösta för det .
Ansvaret för dessa bilar ligger hos tillverkaren .
Det är tillverkaren som måste sörja för infrastrukturen och stå för en rimlig del av skrotningskostnaderna .
Den gemensamma ståndpunkten utesluter inte möjligheten att staten skulle kunna ge bidrag .
Den gemensamma ståndpunkten är en rimlig kompromiss .
En del av dagens ändringsförslag är fullständigt orimliga då de helt och hållet fråntar biltillverkaren ansvaret för att betala en liten del , om ens någon , av skrotningskostnaden för bilar i användning .
Jag kan inte acceptera detta och på skattebetalarnas och de europeiska konsumenternas vägnar röstar jag emot dessa ändringsförslag .
Herr talman , mina ärade damer och herrar !
Det råder enighet om att vi måste börja tänka på hur vi i Europa skall handskas ordentligt med gamla bilar , men rådet har i detta fall inte gett något exempel på en meningsfull europeisk miljöpolitik .
Det var blamerande hur det tyska ordförandeskapet behandlade frågan .
Först stämde Trittin , miljöministern , inte av det hela i tillräcklig utsträckning med sina kolleger i kabinettet , därpå kom förbundskansler Schröder likt en elefant i en porslinsbutik och blandade sig utan sakkunskap i förfarandet .
Men inte heller beslutet från det finländska ordförandeskapet i juni var det bästa man kunde uppnå .
Det finns ett par svagheter .
Den största svagheten är som jag ser det att man inte har tagit tillräckligt stor hänsyn till de medelstora företagens situation , men bilindustrin består inte endast av storföretag .
Just på underleverantörsområdet spelar medelstora företag en mycket stor roll , och vi måste ta hänsyn även till de anställdas intressen i dessa små och medelstora företag .
Därmed är det långt mer än två miljoner människor som har sitt arbete på detta område .
Många ändringsförslag från utskottet för miljö , folkhälsa och konsumentfrågor gagnar just de medelstora företagen , liksom också de föreliggande ändringsförslagen från vår grupp till artikel 5 gällande kostnaderna .
Inte heller från miljöpolitisk synpunkt är den gemensamma ståndpunkten någon lysande prestation .
Det saknas blick för de stora sammanhangen , och när kollegan från De gröna säger att det skulle bli första gången som Europaparlamentet försvagade den gemensamma ståndpunkten så är det ingenting man kan påstå , för ur ett miljöpolitiskt perspektiv är det ju föga meningsfullt om vi genom stela , höga återvinningsmål hindrar moderna , energisnåla fordon såsom 3-liters-bilen , där det ju används mycket plast !
Därför måste man stödja ett ändringsförslag som innebär att man åtminstone tolererar undantag om vi har särskilt sparsamma bilar .
Industrins invändningar är säkerligen inte ologiska på detta område .
Plast- och bilindustrins argumentationskraft skulle emellertid tillta även om man inte bara i detta sammanhang skulle engagera sig för en reducering av koldioxid i Europa .
Herr talman !
I dag befinner vi oss verkligen i en ovanlig situation : De som vill försvara miljövärdena ställer sig bakom rådets gemensamma ståndpunkt .
Till skillnad från föregående talare kan jag konstatera att jag verkligen är stolt över att man under det finländska ordförandeskapet kom fram till en gemensam ståndpunkt som försvarar miljövärdena .
Om vi frångår den gemensamma ståndpunkten och strävar efter att dela kostnaderna för återvinning skapar vi kryphål : Vi får inte något vettigt , klart system där ansvarsförhållandena är i sin ordning .
Därför är det enligt min mening tillverkaren som skall bära huvudansvaret .
Det är bara så vi kan lösa problemet på ett tillräckligt bra sätt och även ta hänsyn till att tillverkarna uppmuntras att tillverka sådana fordon som i framtiden kan återvinnas till så låga kostnader som möjligt .
Herr talman !
Det finns två principiella frågor i rådets förslag till direktiv .
Den ena rör producentens oinskränkta ansvar att återta uttjänta fordon .
Det riskerar att det skapas en monopolsituation inom demonteringsverksamheten .
Särskilt gäller detta i områden inom EU där avstånden är stora , och där många småföretag är engagerade i demontering .
Jag menar att EG : s direktiv inte får , oavsett vad ärendet gäller , missgynna de små företagen inom unionen .
Producenternas oinskränkta ansvar riskerar även att marknaden för begagnade bildelar försvinner .
En producent har ett större ansvar att sälja nya delar .
Denna handel är viktig , särskilt för dem som samlar på och renoverar äldre fordon .
Denna princip är även tveksam utifrån marknadsekonomiska principer .
Företag skall kunna förändras , säljas och avvecklas .
De skall kunna etablera sig på nya marknader , men även lämna gamla marknader .
Att binda producenter med ett ansvar som kan sträcka sig mycket långt bakåt i tiden stämmer illa med en flexibel och utvecklingsfrämjande marknadsekonomi .
Den andra principen i rådets gemensamma ståndpunkt är inslaget av retroaktivitet i direktivförslaget .
Det strider mot vedertagna ekonomiska och juridiska principer , att retroaktivt ålägga en producent ekonomiskt ansvar för sin vara .
Det ändrar även ägaransvaret retroaktivt .
En konsument kan under åren ha ändrat produkten i flera avseenden .
Alla länder inom EU har i dag lagar som reglerar skrotning av bilar .
De kan vara bättre och de kan vara sämre länderna emellan .
I avvaktan på att detta EG-direktiv får genomslag bör emellertid EU-länderna , var för sig , ansvara för skrotning av fordon på bästa sätt , så att retroaktiviteten i EU-lagstiftningen inte tillämpas .
Detta strider inte mot en finansieringsmodell med fonduppbyggnad .
Herr talman !
Att den åtgärd vi diskuterar är viktig för miljön och industrin är uppenbart och någonting vi alla kan enas om .
Den gemensamma ståndpunkten är en godtagbar men mycket känslig och vansklig kompromiss , så mycket mer eftersom den medför ganska begränsade förbättringar om man inte skall äventyra hela direktivet .
Jag hävdar alltså att parlamentet inte kan utöva tvång och att det vore paradoxalt om det skulle göra det om en linje som innebär en minskning av åtgärdens miljökonsekvenser .
Jag påminner om att biltillverkarna har medgett att de kan leva med direktivet .
Kostnaderna är inte astronomiska : att återvinna en bil kostar mindre än 1 procent av nybilspriset .
Dessutom träder tillverkarnas ekonomiska ansvar inte i kraft förrän år 2006 , när en stor del av dagens fordonspark inte längre finns på marknaden .
För de återstående fordonen kan man också införa en slags ansvarsfördelning , såsom föreslås i Langes ändringsförslag 44 och 45 , de enda jag tycker är förenliga med balansen i den gemensamma ståndpunkten och med de aktuella erfarenheterna i somliga länder , och som därför är värda att stödja .
Herr talman !
Detta är ett ytterst dåligt direktiv .
För det första , som min kollega Bowis har påpekat , är det retroaktivt och därför principiellt felaktigt .
För det andra , det lägger enorma kostnader på den europeiska fordonsindustrin , vilket skulle skada konkurrenskraften och sysselsättningen .
I det här parlamentet diskuterar vi ständigt behovet av att främja sysselsättning och arbetstillfällen i Europa och ändå vidtar vi ständigt åtgärder som kommer att ha ett negativt inflytande på sysselsättningen .
Jag vill påstå att direktivet är dåligt även i ett annat avseende , vilket inte har granskats tillräckligt grundligt i denna debatt .
Det är som mycket annat i europeisk lagstiftning .
Det är alldeles för normativt .
Det cementerar en specifik återvinningsmodell .
Det löpande bandet uppfanns för cirka hundra år sedan , jag tror det var av Henry Ford , och det som vi håller på att göra här övertygar mig om att vi försöker skapa något slags omvänt löpande band i artonhundratalsstil - för att demontera fordon , för att ta isär delarna och försöka återvinna dem .
En sak som vi borde tänka på är att marknaden för återvunna stötfångare i plast är mycket osäker .
Plastindustrin vill för det mesta inte ta tillbaka dessa delar och kan av ekonomiska skäl inte heller göra detta .
Det finns redan en mycket framgångsrik industri som skrotar bilar , återvinner metaller och återvinner energi genom förbränning av icke-metalldelar .
Detta är ett ur miljösynpunkt mycket rimligt tillvägagångssätt .
Miljömässigt sett är det lika bra att bränna gammal plast som att bränna ny olja för energiåtervinning .
Denna bilskrotningsmetod medför inga kostnader och skulle sålunda eliminera hela frågan om vem som betalar , eftersom den " döda " bilen i själva verket har ett lågt värde då den kommer in i återanvändnings- och återvinningsprocessen .
Jag motsätter mig detta direktiv eftersom det är för normativt , det tar ingen hänsyn till vad som för tillfället i själva verket pågår på bilåtervinningsmarknaden , och det cementerar metoder som inte nödvändigtvis är de bästa ur miljösynpunkt och säkerligen är mycket skadliga ekonomiskt sett .
Herr talman , kolleger !
Den gemensamma ståndpunkten är bra , men det är parlamentets uppgift att ytterligare förbättra den gemensamma ståndpunkten om uttjänta fordon .
Den socialdemokratiska gruppen har under de senaste dagarna kommit med några viktiga förslag till förbättring .
Jag skulle framför allt vilja göra er uppmärksamma på ändringsförslag 45 .
Där väljer vi att lägga kostnaderna för demontering och återvinning hos producenterna , i alla fall för nya bilar .
I samband med konstruktion och produktion kommer man därigenom att ta hänsyn till återvinning .
För de bilar som nu är i trafik är det rimligt att dela kostnaderna , till exempel genom att inrätta en fond som i Nederländerna .
I den gemensamma ståndpunkten står det att producenterna inte bara skall stå för kostnaderna , utan att de också måste ta tillbaka de uttjänta bilarna .
Det är enligt min uppfattning ett mycket stort problem .
Jag pläderar för att inte låta just biltillverkarna organisera skrotning och återvinning , för det skulle leda till att tillverkarna får ett för stort grepp om marknaden för begagnade delar .
De kan då själva bestämma priserna .
Var och en som någon gång har kört en gammal bil vet att detta är till nackdel för konsumenten och för den som gillar att meka .
Den europeiska konsumentorganisationen , som bett oss att stödja den gemensamma ståndpunkten på den punkten , lämnar enligt min mening konsumenten i sticket .
Ett andra argument för att hålla bilskrotningen borta från tillverkarnas händer är transportkostnaderna .
Om alla biltillverkare kommer att inrätta sina egna skrotningsföretag kommer det att göra det nödvändigt att bogsera bilvrak över långa avstånd .
Det är både miljöovänligt och dyrt .
Inte heller detta har konsumenten någon nytta av .
Därför skulle jag gärna se att ni stöder ändringsförslag 45 .
Herr talman , fru kommissionär !
Jag har återigen begärt ordet för att få säga ytterligare ett par meningar efter den här debatten .
Kära kolleger !
Den som reser till Nederländerna kan konstatera att sista ägaren alltid kan lämna ifrån sig sin bil kostnadsfritt i Nederländerna .
Där kan man konstatera att dessa uttjänta bilar tas om hand på ett meningsfullt sätt , att nya avfallsströmmar har gjorts tillgängliga för att återvinna materialet , att 85 procent av en bils vikt återvinns , att 92 procent av alla bilar återvinns i Nederländerna .
Det finansieras via en fond som nybilsköparna betalar in till .
Fru Breyer , är det ekologiskt förkastligt att så sker ?
Jag svarar nej .
I Nederländerna finns det en förebildlig modell där avfallet efter bilar tas om hand på samma sätt som direktivet föreskriver , och frågan om huruvida det är nybilsköparen som skall betala eller tillverkaren av de gamla fordonen som nu är i trafik har ingenting , över huvud taget ingenting med ekologi att göra utan är en ren fråga om konkurrens !
( Applåder ) Om en europeisk tillverkare skall behöva betala 250 miljoner euro eller en koreansk kanske 2 miljoner euro , det är vad frågan gäller , och precis som människorna som bygger bilar här i Europa är jag för att konkurrensen inte skall gestaltas ojämnt , utan i miljöskyddets anda vill jag att befria sista ägaren från kostnaderna , vilket finansieras genom en fond , och för den nya bilen vill jag naturligtvis att tillverkaransvaret skall gälla , eftersom denne då får bära ansvaret för att tillverka återvinningsvänliga bilar !
( Applåder från PSE-gruppen ) Herr talman !
Det förslag som vi diskuterar innehåller ett mycket stort antal positiva punkter , företrädesvis inriktade på att förebygga avfall , återanvändning , återvinning och recirkulation av delar , återvinning av material och så vidare .
Jag tror att vi har lämnat ifrån oss ett bra förslag .
Diskussionen handlar företrädesvis om ifall konstruktören , den slutliga försäljaren eller någon annan måste ta tillbaka bilvraket gratis eller inte .
Jag skulle bara vilja ta mitt eget land som exempel för att förklara hur det fungerar där utan några problem .
Vi har nått en överenskommelse med alla dem som berörs av denna fråga , det vill säga bilkonstruktörerna , de som handlar med begagnade bilar , bilindustrins samarbetsorganisation , behandlingsanläggningarna för metall , sönderdelningsanläggningarna och staten .
Det finns ett miljöpolicyavtal som undertecknats på frivillig väg .
Bilindustrin , och Belgien är ett land med en mycket stor bilproduktion , har inte ställt till med något som helst problem i samband med detta .
Våra medborgare kan lämna in sin bil gratis till den slutliga försäljaren .
Tvärt emot vad som sägs här , om att detta skulle vara till nackdel för sysselsättningen , har vi kunnat konstatera hur en rad småföretag helhjärtat tagit sig an återvinningen av materialet , och att de gör det på ett mycket bra sätt .
Vissa företag har blivit spetsföretag eftersom de lyckats återvinna vissa material , till och med material som ännu inte är upptagna i direktivet .
Det innebär således att vi här utvecklar en ny sektor , ny sysselsättning och gör miljön en stor tjänst .
Jag är för gratis inlämning .
Det har lyckats hos oss .
Varför skulle det inte kunna lyckas någon annanstans ? .
Herr talman , ärade parlamentsledamöter !
Tack för en intressant debatt med många viktiga argument som har framförts .
Vill ni vara snälla att stå ut med mig under att par minuter .
Tillåt mig att kort redogöra för några av de utgångspunkter och principer som ligger bakom detta direktiv .
Låt mig också börja med att kommentera och svara på ett par av de viktigaste argumenten i denna debatt .
För det första tror jag att vi skall upprepa några grundläggande fakta som redan Florenz och andra har nämnt .
Det vi diskuterar här är det faktum att närmare tio miljoner bilar skrotas varje år i Europeiska unionen , att det utgör ungefär lika många miljoner ton avfall .
Det vill säga närmare tio miljoner ton avfall skapas av dessa bilar , och ungefär 7 procent av dessa lämnas i naturen .
De utgör dessutom miljöfarliga ämnen av värsta slag .
Ungefär 10 procent av produktionen av bly återfinns i bilar , men också kadmium , krom , kvicksilver och andra mycket farliga ämnen .
Detta känner ni redan till , men jag vill ändå upprepa det också för dem som lyssnar .
Detta är en av de snabbast växande avfallsströmmarna som vi har i Europa .
Vi vet att avfallet finns där , vi vet hur vi skall handskas med det , och det finns ingen ursäkt för att undvika att handla .
Det finns tre syften med detta direktiv : För det första vill vi få bort användningen av giftiga tungmetaller från tillverkningen av nya bilar .
Vi vill för det andra slå fast tillverkaransvaret .
Vi kan inte längre ta hand om saker i slutet av en produkts livscykel , utan vi skall undvika att skapa så mycket av avfall .
Vi skall se till att återvinna så mycket som möjligt av en produkts olika innehåll .
För det tredje vill vi nå återvinningsmål som är preciserade i detta direktiv .
Det är de tre viktigaste syftena med direktivet .
Det beror ju på att det är ett slöseri med resurser att vi inte ser till att materialet som finns i bilar återvinns .
Det är framför allt producentens resurser som vi slösar med om vi inte tar itu med en bils livscykel .
Två viktiga frågor har kommit upp här - ja , det finns fler , men jag vill nämna två av de viktigaste .
För det första : Vem skall betala ?
Den andra frågan är : Försämrar vi europeisk bilindustris konkurrenskraft med detta förslag ?
Den första frågan gäller alltså vem som skall betala .
I direktivet framgår det att kostnaden skall bäras huvudsakligen av producenten i enlighet med de principer som vi har i EU : s fördrag om producentansvar samt att förorenaren skall betala .
Det är dock klart att denna kostnad kommer att bäras gemensamt av producenter och konsumenter .
Vi har räknat ut att kostnaden för att återvinna bilar inte utgör mer än en procent av priset för en ny bil .
Tror vi då att kostnaden försvinner , om vi inte skulle anta detta direktiv ?
Nej , det är klart att vi alla kommer att få bära kostnaden för att miljön förstörs , men det blir mycket dyrare .
Dessutom kommer kostnaden längre fram .
Kostnaden försvinner alltså inte , men nu tydliggör vi vems ansvaret är och hur kostnaden skall fördelas .
Talar vi då om en bilindustri i kris ?
Är det en vinstsvag industri som vi diskuterar och som vi verkligen måste hjälpa genom att inte lägga på fler pålagor ?
Är det så att bilindustrin absolut inte har råd ?
Är det så att motiven i själva verket är att försämra europeisk bilindustris konkurrenskraft ?
Nej , naturligtvis inte !
Det är alldeles tvärtom !
Tror ni att konsumenternas krav på miljövänliga bilar och bränslesnålare bilar kommer att minska i framtiden ?
Vad tror ni att barn och barnbarn kommer att ställa för krav på bilar , eller att lagstiftarna i framtiden kommer att ställa för krav på bilar ?
Naturligtvis att de skall vara miljövänliga , att de skall kunna återvinnas , att de skall vara bränslesnåla , att de inte skall förorena vår miljö !
Det är ju bara på detta sätt som vi kan skapa en framtid för bilindustrin .
Vi måste skapa drivkrafter som är sunda , som ser till att vi tar hand om avfallet , att vi återvinner materialet , att vi kan konkurrera med miljövänliga och bränslesnåla bilar .
Det faktum att vi har en europeisk bilindustri som redan är långt framme kompenserar mer än väl att det faktiskt finns fler bilar som de måste ta ansvar för , som rullar i Europa .
Detta är ingen oöverstiglig kostnad eller oöverstiglig uppgift .
Om vi skapar sådana drivkrafter kommer - det är jag helt säker på - marknadskrafterna och de kommersiella intressena i bilindustrin att se till att det växer fram system för att ta hand om både det ena och det andra .
Det kommer att bli allt från försäkringar till bra och vettiga skrotningssystem och återvinningssystem .
Det kommer industrin själv att se till att det uppstår i Europa .
Detta är ingen oöverstiglig kostnad för europeisk bilindustrin .
Det kommer i stället att hjälpa industrin att vara i fronten när det gäller att producera miljövänliga och bränslesnålare bilar så småningom .
Detta måste vi göra för miljöns skull .
Kostnaderna försvinner inte , avfallet försvinner inte .
Annars måste vi alla som skattebetalare eller samhällsmedborgare betala notan ; dessutom blir det dyrare om vi gör det längre fram , ju längre vi väntar .
Detta skulle jag vilja säga inledningsvis .
Jag vill också kommentera frågan om det är retroaktiv lagstiftning .
Om vi räknar med att en bil i genomsnitt lever elva år , menar parlamentarikerna , eller menar någon , att vi skulle vänta elva år framåt i tiden innan vi tar itu med detta problem ?
Menar ni att vi när vi lagstiftar om kemikalier skulle säga att vi inte låtsas om de kemikalier som redan finns på marknaden , och att vi bara lagstiftar för det som skall tillverkas längre fram i tiden ?
Det är klart att vi måste se på det problem som just nu finns där och den utmaning som den existerande bilparken utgör .
Det är fortfarande inget oöverstigligt problem .
Vi kan ta hand om det .
Vi har redan en infrastruktur .
Vi har det som vi behöver för att ta hand om uttjänta bilar .
Jag hoppas naturligtvis att resultatet av omröstningen skall bli bra i dag .
Jag vill också , om jag inte redan har gjort det , tacka Karl-Heinz Florenz för det hårda arbete som han har lagt ned i miljöutskottet på detta förslag .
Det är faktiskt i många avseenden banbrytande vad gäller återanvändning och producentansvar .
Jag tror att det kommer att få mycket positiva och märkbara effekter på miljön .
Vi kan inte fortsätta att blunda för det .
Vi har som sagt både kunskaperna och tillgångar för att klara av detta .
Efter den första behandlingen i Europaparlamentet 1999 hamnade kommissionens förslag i en besvärlig politisk situation i rådet .
Vi fick emellertid en väl avvägd gemensam ståndpunkt i juli under det finländska ordförandeskapet .
Nu måste vi se till att denna lagstiftningsprocess avslutas på ett framgångsrikt sätt .
Det har lagts fram sammanlagt 48 ändringsförslag .
Kommissionen kan anta 10 ändringsförslag helt och hållet .
Tre ändringsförslag kan godtas delvis , och ett kan godtas i princip .
Vissa ändringsförslag rör förbättringar av kommissionens förslag som vi godtog redan vid den första behandlingen , eller återinför i direktivet sådana delar av det ursprungliga förslaget som rådet har tagit bort .
Detta gäller ändringsförslag 5 , utom första delen , 8 , 9 , första delen , 10 , 12 , tredje delen , 15 , 16 , 20 , 22 , 24 och 25 .
Dessa ändringsförslag kan alla godtas .
Ändringsförslag 6 och 21 är nya ; kommissionen kan godta dem .
Kommissionen kan också godta ändringsförslag 26 med vissa redaktionella ändringar .
Jag vill betona att ett antal av de övriga ändringsförslagen som rör förslagets grundläggande komponenter innebär en avsevärd urvattning av den miljöskyddsnivå som är syftet med den gemensamma ståndpunkten .
De kan därför inte godtas .
Parlamentet har av tradition starkt bidragit till att stärka miljölagstiftningen i Europa .
Det skulle förvåna mig och göra mig nedstämd om så inte blev fallet i dag .
Jag är mycket bekymrad över vissa ändringsförslag från parlamentet som ifrågasätter det här förslagets absoluta grundpelare .
Det rör t.ex. utfasning av tungmetaller , tillverkaransvaret och återvinningskravet .
Jag vill bemöta dessa ändringsförslag gruppvis .
Ändringsförslagen 4 , 11 , 12 , 13 , 28 , 30 , 32 , 37 , 42 och 48 gäller utfasningen av tungmetaller .
Ändringsförslag 12 innebär att bestämmelsens ikraftträdande försenas med minst 10 år .
Ändringsförslagen 13 , 28 , 32 , 37 , 42 och 48 innebär att onödiga villkor och undantag införs .
Det skulle innebära att processen med att ersätta de skadliga ämnena kommer att gå långsammare .
Ändringsförslagen 4 , 11 och 30 innebär att tungmetaller måste avskiljas från avfallet före återvinning .
Kommissionen anser att den utfasning som föreslås i den gemensamma ståndpunkten är lättare att tillämpa ur teknisk synvinkel .
Ändringsförslagen 17 , 18 , 27 , 34 , 36 , 38 , 44 och 45 gäller tillverkaransvaret .
Den kompromiss som rådet har kommit fram till är rättvis men skör .
Kommissionen anser inte att ändringsförslagen skulle förbättra balansen utan att samtidigt skapa spänningar .
Jag beklagar den förvirring som uppstod nyligen genom att interna dokument från kommissionen användes på fel sätt , vilket skapade ovisshet om kommissionens inställning i frågan .
Jag vill betona att kommissionen redan 1997 föreslog en särskild klausul om tillverkaransvar , och att kommissionen helt stöder den gemensamma ståndpunkten .
Det lägger inte oproportionerliga kostnader på tillverkarna , långt därifrån .
Ändringsförslagen 39 , 40 , 46 och 47 gäller kvantifierade mål .
Den höga skyddsnivå som den gemensamma ståndpunkten syftar till skulle urholkas mycket om återvinningsmålet för 2006 tas bort .
Dessa ändringsförslag skulle också göra målen besvärliga att handskas med och svåra att övervaka .
Låt mig dessutom kommentera - lyssna noga på vad jag säger nu , eftersom jag har hört detta upprepas i debatten - frågan om veteran- och hobbybilar som nämns i ändringsförslagen 3 , 7 , 9 , andra delen , och 35 .
Sådana fordon omfattas inte av definitionen om avfall och omfattas därför inte av direktivet .
Så vad som än har påståtts här omfattas inte veteranbilar och motorcyklar av direktivet .
Vi anser inte att ändringsförslagen 2 och 14 tillför direktivet något .
Ändringsförslag 23 innebär att kommissionen måste anta kvalitetsnormer för återanvändbara komponenter .
Detta omfattas inte av direktivet .
Det skulle därför krävas ett ad hoc-direktiv från Europaparlamentet och rådet .
Ändringsförslagen 29 , 31 och 41 urvattnar demonteringskraven .
Särskilt ändringsförslagen 31 och 41 riskerar att urholka möjligheterna att återvinna plast , däck och glas .
Kommissionen kan slutligen inte godta ändringsförslagen 1 och 33 av skäl som har med den rättsliga klarheten att göra samt ändringsförslag 19 som kommissionen anser vara onödigt på detta stadium .
Ändringsförslag 43 hör vidare inte hemma i direktivets tillämpningsområde .
Tack så mycket , fru kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer härefter att äga rum .
 
OMRÖSTNING .
( EN ) Fru talman !
Som ni vet är orsaken till att vi röstar om det här betänkandet i dag och inte i förra veckan de talrika översättningsfelen , särskilt i den franska versionen .
Ni har fått en klagoskrivelse av mig angående antalet felaktigheter i detta betänkande samt i andra betänkanden som jag har haft att göra med på sista tiden .
Ett fel som ännu inte har rättats till finns i ändringsförslag 4 .
I den engelska versionen avser vi farmakologiska och vetenskapliga organisationer .
I den franska versionen står det " entreprises pharmaceutiques et organisations scientifiques " .
Kan ni vänligen se till att de fransktalande parlamentsledamöterna får veta att ordet entreprises inte är korrekt .
Det skall inte finnas med i ändringsförslaget .
Och jag ber er igen , fru talman , att se över standarden på de översättningar vi för närvarande får ta emot .
Fru McNally !
Generellt sett är jag själv också bekymrad över att översättningarna ställer till med allt fler problem .
Jag skall höra med enheterna om hur vi skall kunna lösa detta .
( Parlamentet antog resolutionen . )
Betänkande ( A5-0011 / 2000 ) av Langen för Europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets beslut om ett flerårigt program för främjande av förnybara energikällor inom gemenskapen ( 1998-2002 ) - Altener ( C5-0333 / 1999 - 1997 / 0370 ( COD ) ) ( Parlamentet godkände det gemensamma utkastet . )
Betänkande ( A5-0010 / 2000 ) av Ahern för Europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets beslut om antagande av ett flerårigt program för att främja en effektiv energianvändning ( 1998-2002 ) - Save ( C5-0334 / 1999 - 1997 / 0371 ( COD ) ) ( Parlamentet godkände det gemensamma utkastet . )
Betänkande ( A5-0009 / 2000 ) av Graca Moura för Europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets beslut om att inrätta ett enhetligt instrument för finansiering och programplanering för kulturellt samarbete ( Kultur 2000-programmet ) ( C5-0327 / 1999 - 1998 / 0169 ( COD ) ) ( Parlamentet godkände det gemensamma utkastet . )
Andrabehandlingsrekommendation ( A5-0006 / 2000 ) för utskottet för miljö , folkhälsa och konsumentfrågor om rådets gemensamma ståndpunkt ( 8095 / 1 / 1999 - C5-0180 / 1999 - 1997 / 0194 ( COD ) ) inför antagandet av Europaparlamentets och rådets direktiv om uttjänta fordon ( föredragande : Florenz ) ( Talmannen förklarade den gemensamma ståndpunkten godkänd ( efter dessa ändringar ) . )
Betänkande ( A5-0007 / 2000 ) av Berger för utskottet för rättsliga frågor och den inre marknaden om förslaget till Europaparlamentets och rådets direktiv om utstationering av arbetstagare från tredje land i samband med tillhandahållande av tjänster över gränserna ( KOM ( 1999 ) 0003 - C5-0095 / 1999 - 1999 / 0012 ( COD ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Betänkande ( A5-0012 / 2000 ) av Berger för utskottet för rättsliga frågor och den inre marknaden om förslaget till rådets direktiv om en utvidgning av friheten att tillhandahålla tjänster över gränserna till att även omfatta tredjelandsmedborgare som har etablerat sig inom gemenskapen ( KOM ( 1999 ) 0003 - C5-0050 / 2000 - 1999 / 0013 ( CNS ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Betänkande ( A5-0003 / 2000 ) av Marinho för utskottet för rättsliga frågor och den inre marknaden om I. förslaget till rådets beslut om ändring av beslut 88 / 591 / EKSG , EEG , Euratom om upprättandet av Europeiska gemenskapernas förstainstansrätt ( 5713 / 1999 - C5-0020 / 1999 - 1999 / 0803 ( CNS ) ) och II. förslaget till rådets beslut om ändring av beslut 88 / 591 / EKSG , EEG , Euratom om upprättandet av Europeiska gemenskapernas förstainstansrätt ( 9614 / 1999 - C5-0167 / 1999 - 1999 / 0805 ( CNS ) ) ( Genom på varandra följande omröstningar antog parlamentet de två lagstiftningsresolutionerna . )
Betänkande ( A5-0022 / 2000 ) av Brok för utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik om förslaget till rådets beslut om exceptionellt finansiellt stöd till Kosovo ( KOM ( 99 ) 0598 - C5-0045 / 2000 - 1999 / 0240 ( CNS ) ) Fru talman !
Jag skulle bara vilja påpeka att enligt förfarandet medges inte varken att man framlägger eller följaktligen röstar om ändringsförslag i utskottet .
Jag vet inte om detta är enligt reglerna och därför uppmanar jag er att kontrollera om det förfarande som följdes innan denna åtgärd kom till kammaren var korrekt .
Jag noterar det ni just sade , herr Speroni .
( Parlamentet antog lagstiftningsresolutionen . )
Betänkande ( A5-0018 / 2000 ) av Dimitrakopoulos och Leinen för utskottet för konstitutionella frågor om sammankallandet av regeringskonferensen ( 14094 / 1999 - C5-0341 / 1999 - 1999 / 0825 ( CNS ) ) ( Parlamentet antog resolutionen . )
Gemensamt resolutionsförslag om förhandlingarna om regeringsbildningen i Österrike .
Fru talman !
Även på detta område har vi som vanligt ett antal översättningsproblem .
Som utgångspunkt gäller den engelska versionen .
För att ge er ett exempel har det fallit bort något i såväl den nederländska som i den tyska versionen vid punkt 4 liksom vid punkt 5 , och jag citerar de fyra orden på engelska : " in so far as " .
Jag skulle därför vilja be er att använda den engelska versionen som utgångspunkt .
Tack , herr van Velzen .
Jag säger samma sak till er som jag sade till McNally för en stund sedan .
Jag är mycket bekymrad över de översättningsproblem som blir allt vanligare , och jag kan försäkra er att vi kommer att se på detta mycket , mycket allvarligt .
Under alla omständigheter är det givetvis originalversionen som är den gällande .
Fru talman !
Europeiska socialdemokratiska partiets grupp föreslår följande muntliga ändringsförslag .
Jag läser det på engelska eftersom det är resolutionens originalspråk .
" Fördömer Haider för hans förolämpningar mot vissa EU-medlemsländer och deras ledare under de senaste dagarna i uttalanden , som utrikesminister Schüssel har underlåtit att fördöma . "
( Fler än tolv ledamöter reste sig . )
( Parlamentet antog resolutionen . )
Röstförklaringar- Betänkande ( A5-0082 / 1999 ) av McNally .
( FR ) Jag gläder mig åt detta utmärkta betänkande om meddelandet " Kvinnor och vetenskap " !
I detta dokument föreslår kommissionen att vi skall stimulera debatten i syfte att främja kvinnors ökat deltagande i den europeiska forskningen .
Det är ett mål som förtjänar allt vårt stöd .
Utgifterna för forskning och teknik utgör en ansenlig del av Europeiska unionens budget , efter jordbruket och strukturfonderna .
De olika ramprogrammen har inte endast möjliggjort vetenskapliga arbeten av hög kvalitet , utan också ett nydanande samarbete mellan forskare från olika medlemsstater .
Samtidigt finns det få kvinnor inom de vetenskapliga disciplinerna , trots att de uppnår mycket goda resultat under sina studier .
Kvinnornas underrepresentation får inte fortgå .
Därför välkomnar jag med nöje Europeiska kommissionens förslag .
Syftet med detta dokument är en koncentration på åtgärder att vidta på gemenskapsnivå , och mera särskilt via det femte ramprogrammet för forskning och teknisk utveckling , något jag självklart stöder .
Under de kommande åren gäller det att öka kvinnors deltagande , på ett sådant sätt att 40 procent av dem som får Marie Curie-stipendier , deltar i de rådgivande församlingarna och utvärderingspanelerna för hela det femte FoU-ramprogrammet skall vara kvinnor .
För det ändamålet krävs en stimulans av debatten och erfarenhetsutbytet mellan medlemsstaterna , en samordningsstruktur för inrättandet av ett övervakningssystem inom det femte ramprogrammet , kallat " Kvinnor och vetenskap " , vilket bl.a. skall sörja för insamling och spridning av statistik som samlats in under genomförandet av det femte ramprogrammet och som visar hur stor andel kvinnor som har deltagit i forskningsaktiviteterna .
I likhet med föredraganden anser jag att det fordras studier för att analysera orsakerna till skillnaden mellan det antal kvinnor som tar en naturvetenskaplig examen och det antal kvinnor som lyckas få en anställning på det området .
En bättre analys av de hinder som kvinnor stöter på gör att vi kan utveckla en strategi för att undanröja dessa hinder .
Vi måste mobilisera de många nätverken med kvinnliga forskare och få deras hjälp för att formulera en gemensam forskningspolitik .
Europaparlamentet kommer även i fortsättningen att uppmärksamt följa genomförandet av det femte ramprogrammet för FoU , när det gäller främjandet av kvinnor , samt utformningen av idéer till riktlinjer för det femte ramprogrammet .
I fråga om vetenskap , forskning och Europeiska unionens alla övriga politikområden , bör vi integrera genusdimensionen för att sätta stopp för den strukturella diskriminering som hindrar kvinnorna från att konkurrera med lika förutsättningar på arbetsmarknaden . .
( FR ) I sitt meddelande om " Kvinnor och vetenskap " framför Europeiska kommissionen sina goda avsikter att berika den europeiska forskningen genom att mobilisera kvinnorna .
Det är mycket bra och vi gläder oss åt det .
Det finns faktiskt alltför få kvinnor som deltar i forskningsarbeten inom Europeiska unionen .
Vi vet att det enda vi kan göra för att förändra denna situation med underrepresentation av kvinnor inom det vetenskapliga området är att utveckla en utbildningspolitisk inriktning som systematiskt uppmuntrar en diversifiering av unga flickors yrkesval , och då de tagit sin examen vidta positiva åtgärder i arbetslivet .
Men uppenbarligen har vissa kolleger tagit till brösttoner , med tanke på en punkt i betänkandet från utskottet för kvinnors rättigheter och jämställdhetsfrågor som bidrar till förvirring .
En del tolkar den som en kvot , vilken skulle kräva 40 procent kvinnor inom den europeiska forskningen .
Men så förhåller det sig givetvis inte , eftersom en sådan kvot skulle vara orealistisk .
I betänkandet nämns för övrigt inte när en sådan kvot är tänkt att uppnås .
För att skapa lugn och försäkra kollegerna har jag ingivit ett ändringsförslag till resolutionen , där vi helt enkelt noterar att kommissionen i sitt meddelande åtar sig att göra stora insatser för att öka kvinnors deltagande i gemenskapens forskningsprogram , vilket trots allt är hedervärt .
Och varför inte notera att kommissionen skriftligen har meddelat att den anser 40 procent vara ett mycket viktigt mål för kvinnors deltagande på alla nivåer i genomförandet och förvaltningen av forskningsprogrammen .
Detta är inte en kvot !
Det är en mycket välgrundad avsiktsförklaring från kommissionens sida , i den mån det gäller dess egna och inte medlemsstaternas program .
Staterna borde dock komma på den goda idén att för en gångs skull följa kommissionens goda exempel och sätta in lika stora insatser inom ramen för sina egna forskningsprogram .
Men förutsättningen är givetvis att man inser det ! .
( FR ) Det är lyckosamt att det fanns ett så stort samförstånd i debatten om McNallys betänkande , som syftar till att utöka och underlätta kvinnors deltagande i yrken inom området för forskning och vetenskap .
I den här frågan vore det önskvärt att begreppet lika möjligheter får ett bättre genomslag i vardagen , och jag kan endast glädjas åt genomförandet av en politik som bidrar till att kvinnors legitima strävanden tillmötesgås : att få lika tillträde till vetenskapliga studier , att nå ansvarsposter som verkligen står i relation till deras resultat och förmåga , att se snabbt genomförda följdåtgärder som gör att de kan förena familje- och yrkeslivet .
Detta är en nödvändig realistisk och pragmatisk politik , vars syfte är att avskaffa konkreta hinder som har konstaterats vara obestridliga orsaker till denna ojämlikhet .
Men enligt vår mening måste den absolut ta avstamp i begreppet komplementaritet , vilket är det enda som kan rättfärdiga en viljestark politik i frågan .
Det är genom att respektera dessa värden , som verkligen innefattar en respekt för skillnader , och inte genom att luta sig mot ett påstående om en jämlikhet mellan könen - som i sig bär på motsägelser - som vårt reflektionsarbete och åtgärder måste koncentreras på i framtiden .
Det finns i alla fall ingenting som motiverar att man gör det enkelt för sig och bedriver en kvantitativ politik , dvs. att införa kvoter .
Det skulle strida mot det medborgarskapsbegrepp som ledamöterna i UEN-gruppen är särskilt måna om , och det skulle förmodligen få konsekvenser som står i motsats till dem som tycks eftersträvas i McNallybetänkandet , nämligen att kvinnor skall delta i yrken på området för vetenskap och forskning i proportion till deras värde .
Genom att kvinnorna får tillfälle att uppvisa sina verkliga förtjänster och så långt det är möjligt undanröja de hinder som är förknippade med deras särskilda villkor - dock inte inom ramen för en konflikt där de ger intryck av att angripa männens privilegier - kommer de att bevisa intresset av att underlätta utvecklingen av sina yrkeskarriärer , och därmed kommer de att uppnå en förändring av den balans som alltför ofta är till deras nackdel .
Eftersom Europaparlamentet har valt att rösta för en text som uttryckligen vädjar om en kvoteringspolitik , något som jag med stor beslutsamhet försökte kritisera i mitt yttrande , och trots att jag till stor del instämmer i de allmänna riktlinjerna , var jag tvungen att avstå från att rösta om betänkandet av McNally .
Andrabehandlingsrekommendation ( A5-0006 / 2000 ) av Florenz Fru talman , ärade damer och herrar , kära kolleger !
Vi har i dag i en andra behandling röstat om ändringsförslagen till direktivet om uttjänta fordon .
Jag röstade emot hela direktivet , även på grund av att ändringsförslag 34 till artikel 12 och ändringsförslagen till artikel 5.4 inte fann tillräcklig majoritet här i kammaren .
Jag kommer från ett land där 50 procent av EU : s bilpark tillverkas , och det är just det kostnadsfria återtagandet av det gamla bilbeståndet som är kostnadsintensivt och oacceptabelt .
Här kommer enligt min åsikt även arbetsmarknaden att belastas väsentligt genom de kostnader som dessa företag kan vänta .
Detta kan inte vara bra i en europeisk union där vi dagligen funderar kring sysselsättning .
Jag anser att detta är en graverande brist som i princip inte heller passar vårt rättssystem .
Ur denna synvinkel anser jag inte att detta direktiv är godtagbart .
Fru talman !
Jag skulle vilja yttra mig om Florenz betänkande .
Jag tycker att omröstningen har visat att rådets gemensamma ståndpunkt har försvagats men att de stora grupperna här - i synnerhet de tyska företrädarna för de stora grupperna - tack och lov inte lyckades förstöra själva kärnan i direktivet , nämligen producentansvaret .
Tyvärr fick det passera att en effektiv ekologisk politik för avfallsströmmar nu försvagas , nämligen genom den obligatoriska riskbedömningen av ämnen vars hälsovådliga effekter egentligen har varit kända i flera år .
Vi vet att bly , kvicksilver , kadmium och sexvärt krom gömmer stora toxiska faror och hälsorisker och att man genom talrika gemenskapsdirektiv har lyckats minska användningen av detta utan att det har förelegat någon riskanalys .
Här har Europaparlamentet tyvärr böjt sig för industrins intressen .
Jag är likväl mycket glad över att man har inte har lyckats få majoritet för ändringsförslagen från Florenz , Lange och andra , vilka verkligen har försökt baxa ut producentansvaret och överlåta helt åt konsumenterna att stå för kostnaderna för en miljöanpassad hantering av uttjänta fordon .
Jag tycker att det var ett försök som man verkligen borde skämmas över , och jag är glad att det inte lyckades , att man här inte lyckades samla majoritet för det som en stor regering och ledamöterna från en stor medlemsstat försökte sig på , nämligen att på grundval av deras nationella industris intressen dominera Europaparlamentets hållning vid omröstningen .
Fru talman !
Trots att jag tillbringat större delen av mitt liv i snabba bilar håller jag med min kollega Florenz om att man i direktivet om uttjänta fordon måste klargöra att direktivet inte omfattar veteranbilar .
Dessa fina bilar är inte något avfall .
Det var därför jag röstade för ändringsförslagen .
Veteranbilarnas ålder skall inte heller fastställas eftersom det är stora skillnader mellan de nationella bestämmelserna .
På det här sättet kan man bevara historiskt värdefulla fordon för kommande generationer .
Vi får inte heller glömma dem som har veteranbilar som hobby , deras antal överstiger 50 000 bara i Finland .
I stillhet utför de ett mycket värdefullt kulturhistoriskt arbete . .
Processen i parlamentet rörande denna fråga har varit minst sagt förvirrande .
Inför omröstningen i plenum har nya ändringsförslag lagts fram , sådana som redan röstats ned i utskottet .
I den splittrade situation som nu uppstått anser vi därför att rådets skrivningar är de bästa .
Vi behöver ett direktiv på detta område , och därför vill vi också undvika en komplicerad förlikningsprocess .
Direktivet om uttjänta fordon kommer att statuera exempel för kommande lagstiftning .
Det är därför viktigt att producentansvaret är tydligt ; det får inte på något sätt äventyras .
I dag granskar parlamentet för sista gången denna text om så kallade uttjänta fordon och deras öde , dvs. förstörelsen av dem , vilket är en lovvärd avsikt med respekt för vår miljö .
Men det finns två aspekter som man absolut bör beakta i texten .
Först och främst det finansiella ansvaret för denna förstörelse .
Låt oss se till att det inte alltid blir densamme som betalar , dvs. fordonsägaren .
Denne är redan tillräckligt beskattad för sitt fordon som i finansiellt hänseende inte är annat än en bottenlös källa .
Helt nyligen har vi kunnat tala om principen att den som förorenar skall betala , låt oss då tillämpa den förnuftigt och med eftertänksamhet , utan ideologi och utan att ta miste på mål .
Den andra grundläggande punkt som bör återfinnas i denna text , är en uttrycklig föreskrift om att samlarfordon inte skall omfattas av tillämpningsområdet .
På sina håll sägs det att man inte behöver skriva det , eftersom det är uppenbart , men jag är angelägen om att det görs , för vi har allt intresse av att anta tydliga texter .
Låt oss därför rösta igenom dessa ändringsförslag för att bevara bilindustrins juveler .
Dessa antika fordon bär vittne om en kultur och en passion som bör erkännas och respekteras av Europa , i annat fall riskerar vår specifika karaktär att urvattnas .
Det saknas inte exempel bland EU-texterna - i det fallet vet vi att luddighet eller oklarhet inte sällan leder till betydande tvister eller debatter .
Jag skall bara nämna direktiven 79 / 409 och 92 / 43 .
Tydliga texter är en garanti och en rättslig säkerhet för dem som dagligen kommer att tillämpa eller omfattas av dessa texter .
Parlamentsledamöternas kallelse är inte att skapa tvister eller förse domare med rättegångsprocesser , vilka de än är , för då skulle vi inte uppfylla vårt uppdrag .
Vi parlamentariker bör tvärtom anta kristallklara texter för att begränsa tvister . .
( NL ) Att Florenzbetänkandet har gjort så mycket väsen av sig bevisades av den starka lobbymaskin som sattes in , såväl av industrin som av miljörörelsen .
Jag beklagar att konstruktörerna bombarderade Europaparlamentet och rådet med en hel rad argument som antingen inte höll eller som var falska .
Jag vågar säga detta eftersom jag gjorde mig besväret att också ge mig ut på fältet och inhämta upplysningar hos bland annat skrotningsföretag som redan ägnar sig åt återvinning av bildelar med framgång .
De gjorde klart för mig att argumenten om till exempel säkerhetsrisker är struntprat .
Billobbyn lyckades inte i dag , och det är jag glad för .
Direktivet står fortfarande kvar .
Jag räknar med att vi under förlikningen kommer att uppnå ett utmärkt resultat och att ansträngningarna för en bättre miljö vinner över orimliga industriella krav . .
( EN ) Mitt parti har motsatt sig denna åtgärd och de föreslagna ändringsförslagen .
Det finns få saker som är så säkra i livet som skatter , död och miljöförstörelse .
Men det finns inte heller något som är så säkert som att EG : s miljödirektiv har lovvärda syften men i själva verket misslyckas med att uppnå fastställda mål .
När det gäller miljöförstöring liksom synd är vi alla emot den , men för den sakens skull får vi inte tro att varje åtgärd som föreslås mot detta onda med nödvändighet är god .
Faktum är att detta direktiv , liksom så många andra som behandlar miljöfrågor , inte är bra .
Som så ofta är fallet tillför det bara ännu en tung byråkratisk struktur för att kontrollera ett problem , vilket bara tjänar till att skapa flera arbetstillfällen för tjänstemän och kostar motorindustrin och konsumenterna en hel del pengar .
Det enda det inte kommer att göra är att lösa problemet - det är att skjuta myggor med kanoner .
Ingen , inte minst mitt parti , kan vara av någon annan åsikt än att återvinning skall främjas , men det bästa sättet att uppnå detta är att arbeta med marknaden , inte att skapa ett nytt byråkratiskt missfoster .
Ett lämpligare sätt att gynna återvinning är sålunda att lägga skatt på producenter som inte ökar mängden återanvändningsbart material i sina fordon , detta för att med hjälp av skatteincitament och hjälp att rätta sig efter miljökrav uppmuntra privata återvinningsföretag samt skapa incitament för användning av återvunnet material .
Självklart är detta områden där EU inte har någon jurisdiktion och inte heller skall ha någon sådan jurisdiktion .
I avsaknaden av sådan makt , borde man likväl inte försöka ersätta detta med en mindre effektiv åtgärd .
I stället borde man låta medlemsländerna utveckla sina egna system och undvika tendensen att ingripa där detta inte är önskvärt eller gör någon nytta .
Betänkande ( A5-0007 / 2000 ) av Berger Med detta förslag till direktiv vill man fastställa villkoren för utstationering av arbetstagare från tredje land i samband med tillhandahållande av tjänster över gränserna .
Nationaliteter från tredje land med legalt uppehållstillstånd i en medlemsstat åtnjuter inte rätten till fri rörlighet i Europeiska unionen .
Hittills har det varit stränga restriktioner i den fria rörligheten för arbetstagare från länder utanför unionen .
Det är alltså positivt att man underlättar rörligheten för arbetstagarna i Europeiska unionen , även för arbetstagare från tredje land .
Emellertid syftar bara diektivförslaget till att tillåta deras förflyttning till en annan medlemsstat när det är i arbetsgivarens regi , en arbetsgivare som är etablerad i ett land där han också har sin hemvist , men möjligheteten till rörlighet är begränsad till tiden för utstationering , och bara till den medlemsstat där arbetstagaren har blivit utstationerad .
Detta innebär att det främsta syftet med detta förslag inte är att lösa problemet med dessa arbetstagares rörlighet , utan bara att skapa bättre villkor för företagen som tillhandahåller tjänster .
Å andra sidan för att underlätta förfarandena tas det i Bergerbetänkandet upp ändringsförslag som är djupt diskutabla , vilket skapandet av ett gemensamt informationssystem om tillgång till kort EG-kort utgivna av en myndighet i någon av medlemsstaterna är ett exempel på .
Betänkande ( A5-0007 / 2000 ) och ( A5-0012 / 2000 ) av Berger .
( FR ) Det är med största tillfredsställelse som jag välkomnar de två förslag till direktiv som syftar till att underlätta den fria rörligheten för arbetstagare från tredje land och samtidigt det fria tillhandahållandet av tjänster .
Dessa förslag går i huvudsak ut på att införa ett EG-kort för tillhandahållande av tjänster , som i framtiden kommer att ge nära 5 miljoner medborgare från tredje land som vistas legalt i en av Europeiska unionens medlemsstater möjlighet att tillhandahålla tjänster i andra medlemsstater , något som i dag hindras av problem med att få visum och arbetstillstånd .
Det första förslaget i direktivet skall tillåta de företag som är etablerade i en medlemsstat och som har arbetstagare från tredje land att tillfälligt utstationera dessa arbetstagare i en annan medlemsstat för att tillhandahålla tjänster där .
I enlighet med de föreskrivna bestämmelserna skall arbetsgivaren bara behöva göra en förfrågan om ett kort för tillhandahållande av tjänster för varje berörd arbetstagare .
För att kunna få ett sådant kort bör arbetstagaren logiskt sett vistas legalt i en medlemsstat och omfattas av ett socialförsäkringssystem .
Det andra förslaget ger samma rättigheter åt egna företagare från tredje land .
Innehållsmässigt ansluter jag mig till Europeiska kommissionens förslag .
Vissa bestämmelser kan dock skapa förvirring , och därför röstar jag för de ändringsförslag som har ingivits av föredraganden .
De kan bidra till att bestämmelserna tydliggörs och således till att man förekommer alla former av missbruk !
Andra ändringsförslag syftar till att förenkla de administrativa förfarandena , till exempel genom att låta medlemsstaterna utse en myndighet som skall ha ansvaret att utfärda korten .
En sådan ändring verkar nödvändig för att undvika det byråkratiska krångel som alltför ofta bromsar en bra tillämpning av nya bestämmelser .
Därför kan jag bara glädja mig åt att dessa ändrade direktiv har antagits , eftersom vi inte mycket längre kan acceptera att personer som under lång tid har vistats legalt inom Europeiska unionen skall stöta på så många svårigheter .
Det går stick i stäv med den grundläggande princip om icke-diskriminering som är inskriven i unionens grundfördrag .
Betänkande ( A5-0003 / 2000 ) av Marinho Rådets förslag till ändringar har väckt starka reservationer från vår sida .
För hur kan man förklara att det behövs fler domare vid förstainstansrätten , som man vet är överbelastad , och samtidigt föreslå att rättens behörighetsområde skall utökas ?
Den första åtgärdens effekter tillintetgörs de facto av den andra .
Vissa skulle säga att det inte finns något sådant som perfektion , men en kort historisk påminnelse borde göra det lättare för dem att förstå våra förbehåll : Den 1 januari 1995 tog rådet åter upp frågan om ett ökat antal domare i enlighet med artikel 17 i anslutningsfördraget av den 24 juni 1994 .
Redan under förberedelsen av Amsterdamfördraget i maj 1995 oroades förstainstansrätten över det ständigt ökande antalet mål , och insisterade på att det krävs åtgärder , " i annat fall kan rätten snart inte till fullo uppfylla principen om god rättsförvaltning och ombesörja det uppdrag som den har anförtrotts ... omständigheterna är sådana att skyddet av dem som står i kontakt med rättvisan kan äventyras " .
Vad gjorde man då i Amsterdam ?
Ingenting i den riktningen ; tvärtom ökade bördan då gemenskapens rättsliga befogenheter utökades inom områden som tillhör den tredje pelaren .
Ni är dessutom överens om att de texter som kammaren röstar igenom alltid vädjar om en domsrätt för gemenskapen , även när det gäller stadgan om de grundläggande rättigheterna som just nu utarbetas .
Det är ingen lösning att förstainstansrätten får 21 domare i stället för 15 eller att rätten , som nyligen , bereds möjligheten att i vissa ärenden vara domför med en domare , det är helt enkelt illusioner som man motvilligt har gått med på och som utsätter oss för alltför sent påkomna insikter .
Dessa förslag är således inte i nivå med det som står på spel , de är ett uttryck för att man går för snabbt fram genom att på sikt kräva flera hundra domare .
Vi kan inte gå med på det , eftersom tendensen till ett domarnas Europa skadar ett gott utövande av demokratin i våra stater .
Enligt vår mening verkar det vara dags att inleda ett grundläggande reflektionsarbete för att få ordning på gemenskapens rättssystem och garantera en rättskipning med kvalitet .
Den frågan går inte att särskilja från den pågående reflektionen om en normhierarki och en bättre tillämpning av subsidiariteten .
Är inte den kommande regeringskonferensen det bästa tänkbara tillfället ?
Betänkande ( A5-0018 / 2000 ) av Dimitrakopoulos och Leinen .
Den stundande regeringskonferensens viktigaste uppgift är att reformera EU inför mottagandet av de nya medlemsländerna .
Vi stöder därför givetvis att Europaparlamentet nu ger sitt formella klartecken till att regeringskonferensen startar .
Vi anser dock att regeringskonferensen skall begränsas till frågor som är nödvändiga för att utvidgningen skall kunna göras .
Detta hävdade vi också i november 1999 , och vi vill därför hänvisa till vår röstförklaring av den 18 november 1999 . .
( FR ) I den ståndpunkt som Europaparlamentet just har antagit om inledningen av nästa regeringskonferens , vädjar parlamentet om att man bör " inleda en konstitutionell process " .
Denna vilja att kontrollera nationerna med en juridiskt sett högre stående text kommer också till uttryck på de första sammanträdena i den församling som har i uppdrag att utarbeta en så kallad stadga om de grundläggande rättigheterna , men i realiteten en maskerad konstitution .
Den viljan uttrycks också i det osannolika steg som i dag tas i Europaparlamentet : önskan att radera resultatet av de fria valen i Österrike genom att rösta igenom en resolution .
Samma vilja att göra nationerna till vilka underordnade administrativa regioner som helst , framgår också av alla sidorna i kommissionens yttrande inför regeringskonferensen .
Den centrala idén består i att generalisera omröstningarna med kvalificerad majoritet och samtidigt förändra innebörden av denna kvalificerade majoritet , genom att omvandla den till en dubbel enkelmajoritet - staterna och befolkningarna - med syftet att öka kommissionens handlingsutrymme och minska densamma för de stater som är i minoritet .
Fransmännen kommer utan tvekan att vara intresserade av att - så här i förbigående - få veta att kommissionen begär en ändring av artikel 67 i Amsterdamfördraget för att där införa majoritetsomröstningar , samt ett medbeslutande med Europaparlamentet .
Man bör minnas att denna artikel , som handlar om invandringspolitikens överföring till gemenskapspelaren , föreskriver att besluten skall fattas enhälligt i rådet under fem års tid , och att rådet sedan skall bedöma om det eventuellt är lämpligt att ändra på systemet .
I Frankrike , både i nationalförsamlingen och i senaten , kände sig många parlamentsledamöter lugnade när fördraget ratificerades , eftersom man sade att rådet under alla omständigheter kommer att ha frihet att välja och att det därmed skulle kunna bevara enhälligheten .
Men i dag föreslår Barnier - den Europaminister som förberedde Amsterdamfördraget och som under tiden har blivit ledamot av Europeiska kommissionen - att man vid nästa regeringskonferens skall besluta att rådet skall arbeta på de här frågorna med majoritetsbeslut .
Detta är ett exempel på att vi ständigt hamnar i en ond cirkel när vi spelar spelet om den europeiska integration med institutionerna i Bryssel .
Fransmännen måste inse att alla dessa åtgärder inte endast syftar till att deras land skall försvinna såsom ansvarigt beslutscentrum , utan att man också kommer att utnyttja alla medel för att avtvinga dem deras samtycke till detta .
Ger de efter är de förlorade .
För det man håller på att ta bort , det är deras försvarsmedel , ett efter ett . .
( DA ) De danska socialdemokraterna har i dag röstat emot betänkandet om sammankallande av regeringskonferensen .
Det är avgörande för oss att denna regeringskonferens kan avslutas före utgången av år 2000 , så att det inte blir formella förhållanden som röstviktning i ministerrådet och sammansättningen av kommissionen och Europaparlamentet som lägger hinder i vägen för utvidgningen av EU .
Vi var därför också mycket nöjda med de beslut som fattades om detta på toppmötet i Helsingfors i december .
En alltför ambitiös utvidgning av dagordningen vid nuvarande tidpunkt riskerar att försena utvidgningsprocessen .
Detta vill vi inte skall ske - vi har därför röstat emot .
Vi håller emellertid helt med våra kolleger om att det finns behov av öppenhet i samband med regeringskonferensen , så att medborgarna får klart för sig hur arbetet fortskrider . .
Vi är nöjda med att det sattes upp en begränsad dagordning för regeringskonferensen vid mötet i Helsingfors .
Utformningen av det framtida EU bör även eventuella blivande medlemsstater vara med och ha ett inflytande över .
Valet till Europaparlamentet 1999 visade med all tydlighet att medborgarna inte följer med i tankegångarna om ett allt mer Brysselfederalistiskt EU . .
( FR ) När nästa regeringskonferens inleds blir Europeiska unionens metod åter aktuell .
Än en gång kommer stats- och regeringscheferna att skaffa sig ensamrätt till debatten .
Det betyder att femton personer kommer att diskutera och fatta beslut inom lykta dörrar om 350 miljoner människors framtid .
Man kan därför förstå folkens ointresse för ett europeiskt bygge som uppförs bakom ryggen på dem och långt ifrån deras angelägenheter .
Det räcker faktiskt med att titta på regeringskonferensens dagordning : institutionerna , utvidgningen och ett självständigt försvar .
I realiteten handlar det om att förstärka den verkställande makten , att utveckla östländernas införlivande av liberalismen och att driva på en militarisering av Europa , bl.a. genom att utöka försvarsbudgetarna .
Det sociala Europa , något som EU framhåller , har helt enkelt försvunnit från dagordningen .
Allt detta legitimerar bara utvecklingen av motståndsrörelser på Europanivå , rörelser som vill införa en social stadga för att arbetstagarnas viktigaste krav skall harmoniseras ovanifrån .
Därför röstar jag emot betänkandet .
Jag röstade för resolutionen som är positivt till sammankallandet av en regeringskonferens eftersom det befäster det portugisiska ordförandeskapets filosofi , med stöd från en stor majoritet i parlamentet , om att öppna regeringskonferensens dagordning för andra frågor än de som är strikt relaterade till maktbalansen mellan medlemsstaterna , stora och små , så som ursprungligen fastställdes i kallelsen till rådet i Helsingfors .
Tyvärr är de ämnen som tas upp i resolutionerna om de framtida frågorna för en revidering av fördraget om behovet att se över artikel 7 , som handlar om avstängning av en medlemsstat om den på ett allvarligt och återkommande sätt kränker unionens ursprungliga principer i artikel 6 .
Så som visas i den nuvarande krisen med Österrike , har unionen rätt att försvara sig .
Emellertid är de rättsliga mekanismerna som finns i fördraget svaga , och svåra att tillämpa politiskt och rättsligt , de klassificerar inte institutionernas makt och garanterar inte en rättslig behandling av en process av större betydelse vilket just ett fördömande och avstängning av en medlemsstat innebär .
Därför anser jag att denna fråga genast måste föras upp på regeringskonferensens dagordning , och detta motiverar i sig en långtgående revidering .
De frågor , som vi för närvarande anser vara centrala , när det gäller sammankallande av en regeringskonferens för att revidera fördragen är långt viktigare än kontroversen här angående varje dagordnings dimension , när det gäller möjligheten att formulera förslag till nya frågor att ta upp och Europaparlamentets deltagande i den .
De relevanta frågorna , enligt vår mening , handlar om regeringskonferensens möjligheter och syften och de frågor som kommer att debatteras .
Vi tvivlar på möjligheterna eftersom vi har de verkliga målen i sikte , kanske långt ifrån det alltid nämnda anpassningen till den planerade utvidgningen .
Detta syns särskilt i det innehåll som eftersträvas , speciellt inom de områden som ej löstes i Amsterdam - och detta tyder på ett framtida skapande av oacceptabla direktorat - , men också för det som handlar om andra och tredje pelaren , vilka tenderar i en riktning mot en oönskad militarisering av Europeiska unionen .
Det här är några av de främsta skälen till att vi inte stöder inriktningen av detta resolutionsförslag .
Europeiska socialdemokratiska partiets grupp lade ned sina röster vid den senaste omröstningen om betänkandet av Leinen Dimitrakopoulous .
Texten är överambitiös , och Storbritanniens parlamentsledamöter från Labour anser att regeringskonferensen i första hand borde behandla " resterna av Amsterdam " , detta för att förbereda utvidgningen och inte breda ut sig alltför mycket utanför detta .
Det pågår för närvarande en hel del reformarbete , och detta måste för tillfället prioriteras för att möjliggöra en konsolidering och förstärkning av EU : s institutioner .
En utökning av dagordningen och en drastisk revidering av fördragen skulle föra med sig en risk för destabilisering .
Huvudfaktorn i den här texten , såsom ändringsförslaget lyder , är en begäran om att en stadga om grundläggande rättigheter skall införlivas i fördragen .
Enligt vår mening skulle detta medföra en komplicerad lagstiftningsbörda .
En politisk och fastställande stadga , som för medborgarna klargör deras gällande rättigheter , vore att föredra .
Vår prioritering ( dvs . " resterna " ) måste vara : antalet kommissionärer samt deras ansvar röstviktningen i rådet utvidgningen av den inre marknaden inom områden som gynnar Storbritannien och Europa ( men inte fördragsändringar , försvarsfrågor , gränskontroller eller beskattning ) och inslaget av medbeslutande på områden dit den inre marknaden utvidgats Utöver detta befarar vi att " flexibiliteten " eller förslaget om ökat samarbete inte är lämpligt för närvarande .
Amsterdam-bestämmelserna är till stor del oprövade och att skapa ett större utrymme för avhopp skulle försvaga EU i ett skede då man överväger en utvidgning och då ansökande länder uppmanas att anpassa sina lagar till en inre marknad och annan europeisk lagstiftning . .
För att kunna påverka utvecklingen måste Europaparlamentet inta en mer konstruktiv attityd till regeringskonferensens dagordning än som framkommer i denna resolution , vilken i alltför stor utsträckning ägnar sig åt besvikelse och negativism över det beslut som Europeiska rådet fattade i Helsingfors i december 1999 .
Europaparlamentet och dess konstitutionella utskott borde i stället ha preciserat sig och koncentrerat sig på några få punkter utöver rådsbeslutet i Helsingfors och därmed ange vad man anser vara mest angeläget att ta upp till behandling , bland annat frågan om inrättande av en åklagare för brottslighet riktad mot Europeiska unionens institutioner och deras ekonomiska intressen .
Vi svenska kristdemokrater motsätter oss också hot om att försena östutvidgningen av EU som framförts om inte regeringskonferensen utvidgas mycket omfattande utöver vad som blev kvar från förra regeringskonferensen i Amsterdam 1997 . - Den stundande regeringskonferensens viktigaste uppgift är att reformera EU inför mottagandet av de nya medlemsländerna .
Jag stöder därför givetvis att Europaparlamentet nu ger sitt formella klartecken till att regeringskonferensen startar .
Jag anser dock att regeringskonferensen skall begränsas till frågor som är nödvändiga för att utvidgningen skall kunna genomföras .
I övrigt hänvisar jag till min röstförklaring av den 18 november 1999 där jag klargör min inställning gentemot överstatlighet och ett gemensamt försvar .
Gemensam resolution om Österrike Fru talman !
Gruppen Nationernas Europa har inte anslutit sig till PPE-DE- och PSE-gruppens gemensamma resolution om den politiska situationen i Österrike , vilken uppstått till följd av att de konservativa och Jörg Haiders nationalliberaler bildat koalitionsregering .
PPE-DE- och PSE-gruppens resolution applåderar det initiativ som togs av fjorton medlemsstater för att sätta press på Österrike , genom att organisera en sorts diplomatisk bojkott .
Det som chockerar oss mest är att denna gemensamma intervention viftar med fördragets principer som om det någonstans stod skrivet att ett folks fria och demokratiska uttryck kan upphävas av grannländernas stats- och regeringschefer , som för övrigt har aktat sig noga för att samråda med sina respektive folk .
Vilka verbala övertramp Jörg Haider än har gjort , och vi beklagar faktiskt dem , har österrikarna gjort ett demokratiskt val , och det måste vi respektera .
I våra ögon är det uppenbart att vänstern i Europaparlamentet - i samförstånd med den österrikiska vänster som besegrades i striden om väljarna - har iscensatt en ren och skär politisk operation som för tankarna till en olycksbådande epok , men som vi lyckligtvis har lämnat bekom oss .
Även om jämförelsen mellan Haider och Hitler saknar all trovärdighet , har den delvis fyllt sin funktion genom att få vissa PPE-DE-ledamöter att vackla .
Men bortsett från denna politiskt förslagna operation , finns det en sak som majoriteten i Europaparlamentet särskilt fruktar , och det är att ifrågasättandet av vänsterns och högerns sammanboende i Österrike - något som har fördärvat det politiska livet - snart sprider sig till det europeiska systemet med gemensamt styre , ett styre som ger upphov till lika beklagansvärda effekter .
För att undvika ett sådant ifrågasättande är denna majoritet beredd till allt : att sudda ut resultaten av fria val ; att inrätta en tankepolis ; att införa en ny form av totalitarism .
Fru talman !
För ledamöterna från Nationella fronten , Vlaams Blok och den italienska sociala rörelsen vill jag ställa följande fråga : vem är det som drar i trådarna i den förskräckande inblandning i Österrikes inre angelägenheter som Europeiska unionen har hängett sig åt i strid med den allmänna internationella rätten , i strid med fördragen , i strid med moralen ?
Är hysterin spontan ?
Är den en frukt av ren dumhet eller - mera troligt - av en avsiktlig strategi , densamma som brukas överallt annars i världen ?
Vem dikterar sin vilja för de europeiska nationerna och gör anspråk på att förbjuda dem att välja ett eget öde ?
Hemliga nätverk ?
Regeringen i Washington ?
Den i Israel ?
Eller deras socialistiska reservtrupper , som i denna församling har fräckheten att sprida sina värderingar bland oss ?
Vilka är då socialisternas värderingar , de socialister som har nått stora valframgångar under det senaste seklet genom att förespegla de sämst lottade en större social rättvisa , men som i dag inte är mer än ett parti för skyddade tjänstemän , etablerade fackföreningar och statskapitalism ?
Vilka är det belgiska socialistpartiets värderingar , ett parti som går från pedofilskandaler till korruptionsaffärer , till att börja med Vandamaffärerna , såsom Agustaaffären ?
Vilka är värderingarna inom det franska socialistpartiet , som i Urba- , Sages- och Graco-affärerna har övat utpressning mot alla de kommuner som är beroende av socialisterna ?
I François Mitterrands parti , Mitterrand som tilldelades Vichyregimens emblem av Pétain , har de högsta ämbetsmännen just blivit tagna på bar gärning , när de levde gott på att förskingra offentliga medel avsedda till en sjukförsäkring för studenter .
Jag skall inte ta upp det italienska socialistpartiets korruptionsaffärer , för man slår inte på den som redan ligger , och än mindre på den som redan är död .
Jag skall däremot tala om det spanska socialistpartiet , som just har ingått en allians med slaktarna från Albacète som gjorde upp med de baskiska nationalisterna med hjälp av lejda mördare .
Jag kommer att tala om det tyska socialistpartiet , som har för avsikt att undervisa oss om andra världskriget - ett international-socialistiskt parti , precis som dess likar var national-socialistiska , som fortfarande marscherar , Waffen-SS : s parti ...
( Talmannen avbröt talaren . )
Fru talman !
Jag har haft stora svårigheter med denna resolution .
Till slut lade jag av flera orsaker ned min röst .
Jag sympatiserade med EDD-gruppens ändringsförslag , som behandlar förkastandet att EU : s ingriper i bildandet av regeringar i medlemsstaterna , men jag var tvungen att lägga ned min röst , eftersom förslaget precis följde på fördömandet av främlingsfientlighet , rasism etc. och jag tyckte att det kunde misstolkas .
Men jag funderar över hur klokt detta är .
För det första uppstår frågan om bekämpning av intolerans med intolerans och de långsiktiga följderna av detta .
Jag undrar också hur klokt det är av EU att reagera på regeringsbildningen i Österrike och hur detta kommer att påverka den allmänna opinionen där .
För tillfället verkar det som om Haiders parti snarare får mera stöd än mindre från oppositionen i utomstående regeringar .
Till och med USA har nu meddelat att man överväger att bryta de diplomatiska förbindelserna .
Vi undrar om detta inte i själva verket underblåser främlingsfientligheten och gagnar de partier och människor som understöder detta .
Jag tycker verkligen att folk borde vara väldigt försiktiga .
Om man vill bekämpa främlingsfientlighet och rasism , och jag tror att vi måste det , måste vi fokusera på grundorsakerna .
Vi måste iaktta de människor som röstar på dessa partier och förstå varför denna situation uppstår .
Det är ingen situation som de flesta i detta parlament önskar , men vi måste vara försiktiga i vårt val av synsätt , så att vi inte till slut åstadkommer raka motsatsen till det vi försöker uppnå .
Fru talman , kära kolleger !
Jag avvisar varje sorts främlingsfientliga och rasistiska uttalanden , manifestationer eller känslor .
Jag försvarar intensivt de mänskliga rättigheterna och rättsstaten , vilket Europa består av .
Men jag är ändå oense med det befängda agerandet som ordförandeskapet ( tyvärr det portugisiska ordförandeskapet ) har initierat i en verkligt institutionell dumhet för fjorton andra medlemsstaters räkning .
Detta är inte ett sätt att bekämpa extremism på .
Det kan till och med vara ett sätt att spela dem i händerna på ett oöverskådligt sätt .
Den kaskad av förvirrade och förhastade åtgärder som vräkts över Österrike blandar ihop allt på ett oproportionerligt sätt , och det stör många medborgare med god vilja och utgör risker som inte har beaktats .
Det finns en oförenlig motsättning mellan ståndpunkter som tas i de mänskliga rättigheternas och rättsstatens namn , men som , samtidigt förolämpar österrikarna i grundläggande rättigheter och kör över de grundläggande rättigheterna i en rättsstat , i detta fall fördragets bestämmelser .
Vad vill vi när vi inleder en regeringskonferens ?
Ett Europa med 27 länder eller ett Europa med 14 , eller ännu mindre ?
Vi är för Europa , ett Europa som hedrar alla de steg vi har tagit för att komma hit , ett Europa som respekterar fördragen och lagen , ett Europa där Österrike behövs .
Det är viktigt att säga detta !
Fru talman !
Jag är glad och stolt över att detta parlament , med övervägande majoritet , har fördömt bildandet av koalitionen i Österrike med Haiders liberala parti .
Haider har under de senaste åren såväl i ord som handling visat att han förtjänar att utestängas från en vanlig demokratisk dialog .
Han har inte bara beundrat Adolf Hitler , berömt Waffen SS och vägrat fördöma en terroristattack som dödade fyra romer , han har också varit ledamot i det regionala styret i Kärnten .
Han har lett satsningar för att dra in bidrag åt Österrikes slovenska minoritet och stöd åt immigranter .
En del har hävdat att vi inte har rätt att ingripa i österrikisk politik .
De har fel .
Genom Europeiska unionens fördrag är vi förpliktade att skydda grundläggande rättigheter .
En del har hävdat att vi måste acceptera resultaten av demokratiska val .
Men demokratiska val gör inte demokrater av dem som har hotat demokratin .
För dem som hävdade samma sak med avseende på Tyskland under 1930-talet , finns det ett tragiskt minnesmärke i form av Förintelsen - 6 miljoner judars död .
Men vi skall inte döma Haider för hans ambition .
Somliga människor ändrar aldrig åsikt .
De skyldiga är egentligen kristdemokraterna i Österrike som beter sig som syndabockar för att återuppliva det hot mot Europa som vi trodde dog i Berlin 1945 .
Fru talman !
Vi har nyligen antagit en resolution som fördömer Jörg Haiders liberala partis rasistiska och främlingsfientliga förflutna i Österrike .
Detta har gjort det möjligt för våra regeringar att handla genom att bryta de politiska förbindelserna med varje regering som han är medlem i och visar också vårt stöd för anti-rasistiska grupper inom den demokratiska majoriteten av Österrikes folk .
Vi varnar för att den här koalitionen , om den bildas i dag , på ett oacceptabelt sätt legitimerar extremhögern , i direkt motsats till de principer om fred och försoning som för oss samman i denna Europeiska union .
Detta är de värderingar vi önskar se hos dem som vill gå samman med oss .
Europaparlamentet kräver att Europeiska kommissionen är vaksam när det gäller rasistiska aktioner i Österrike och hotar med att utesluta Österrike som medlem ur Europeiska unionen om sådana förekommer .
Jag är stolt över att understödja en sådan resolution .
Trots att vårt förslag om att dra tillbaka alla politiska inbjudningar till österrikiska regeringsföreträdare till Europaparlamentet inte antagits i dag , vill jag meddela att vi kommer att fortsätta med att driva detta förslag för att säkerställa att Europaparlamentet gör allt som står i dess makt för att bekämpa återkomsten av nynazister till regeringar i Europa .
Fru talman !
Jag skall fatta mig mycket kort .
Jag respekterar parlamentets önskan som den har framkommit , men jag måste också säga att folkens rätt till självbestämmande inte kan ifrågasättas ens av Europaparlamentet .
Handlingen är orättvis gentemot våra österrikiska kolleger , både nationella och europeiska parlamentsledamöter , och luktar misstänksamhet och politiska , men också kommersiella , intressen lång väg .
Jag tycker inte att man botar medborgarnas ointresse för Europa med dessa signaler .
Den österrikiska extremhögern har fått en oförtjänt present .
Jag uppskattade de italienska radikalernas ståndpunkt mycket , och det säger jag utan att förglömma de historiska och faktiska skillnaderna mellan italienska och österrikiska liberaler .
Jag har under många år i ord och handling varit engagerad i den antifascistiska kampen , kampen för jämställdhet och kampen mot främlingsfientlighet .
Men det som skett under den senaste tiden , först i samband med det som i verkligheten var problem inom ministerrådet , sedan med ordförande Prodis problem med den österrikiske kommissionären och senast i och med denna resolution , är inte något jag kan ställa upp på .
Jag har inte kunnat rösta för denna resolution , även om jag stöder vissa slutsatser .
Det handlar först och främst om en illavarslande blandning av makt , arrogans och svaghet från den Europeiska unionens sida .
Dessa åtgärder strider inte bara mot fördragen och ger unionens organ mer maktbefogenheter än vad som tillkommer dessa , utan det värsta är att de kommer att motverka sitt eget syfte .
Det kommer inte att försvaga Haider och FPÖ ( Österrikiska liberala partiet ) , det kommer tvärtom att stärka dem .
Vi uppnår det rakt motsatta .
På detta sätt bekämpar man inte rasism och högervridning . .
( DA ) Venstres ledamöter vid Europaparlamentet lägger vikt vid att parlamentet vid antagandet i dag INTE har stött de fjorton statsministrarnas diplomatiska sanktioner mot Österrike .
Därför stödde Venstres ledamöter vid parlamentet det liberala beslutets kraftfulla avståndstagande från varje form av främlingsfientlighet i Österrike och på andra ställen .
Vi fäster avgörande vikt vid att Amsterdamfördragets nya bestämmelser används om detta är nödvändigt , så att ett land som i handling kränker grundläggande medborgerliga rättigheter genom diskriminering e.d. , fråntas rösträtten i EU : s ministerråd ( art .
7 ) . .
( EL ) FPÖ : s deltagande i Österrikes regering innebär en mycket stor fara för Europeiska unionens fortsatta politiska utveckling .
Det rör sig om " ormens ägg " som nu tyvärr åter dyker upp i Europa , starkare än någonsin sedan andra världskriget .
Europaparlamentet och unionens regeringar är skyldiga att politiskt isolera en regering som innehåller anhängare av nazism och främlingsfientlighet .
Europeiska unionen - och samtidigt de båda dominerande politiska riktningarna , socialdemokrater och kristdemokrater - har ett stort ansvar , för det är genom EMU : s dogmatiska och stränga budgetpolitik , nedrustningen av välfärdsstaten och hyllandet av den tygellösa konkurrensen som stora befolkningsgrupper har marginaliserats , och därigenom har högerextremistiska demagoger av Haiders typ fått möjlighet att mobilisera anhängare till sin nynazistiska politik . .
( FR ) Eftersom Europaparlamentets bestämmelser inte tillåter oss att lägga fram en egen resolution för att fördöma Haiders parti , liksom alla partier från vilket europeiskt land som helst som sprider rasistiska , främlingsfientliga och illvilliga tarvligheter mot invandrade arbetstagare , har vi röstat för kompromissresolutionen utan att stämma in i flera bedömningar och ordalag , för att visa vår solidaritet med dem i Österrike som motsätter sig den österrikiska extremhögern och dess demagogi .
Vår röst innebär på intet sätt en garant för de partier som undertecknat kompromissresolutionen , varken för deras nuvarande politik eller deras framtida attityd i händelse av ett ökat hot från extremhögern .
Vissa av dessa partier , som ger sig ut för att vara republikanska och demokratiska , har anammat extremhögerns demagogi - av medbrottslighet eller valtaktiska skäl - om så bara för att - öppet eller på ett hycklande sätt - göra de invandrade arbetstagarna ansvariga för arbetslösheten och försvåra deras liv .
De personer från de undertecknande partierna som leder eller har lett en regering i Europeiska unionens olika länder , har på ett mera allmänt plan en del av ansvaret för extremhögerns nyförvärvade inflytande , eftersom de bedriver en politik som av lojalitet med de stora arbetsgivarnas intressen saknar åtgärder för att bekämpa arbetslösheten och den misär som följer i dess fotspår , och därigenom underblåser extremhögerns främlingsfientliga demagogi . .
( FR ) Den här veckan har Europa utan tvivel gett till sitt första politiska skrik .
Genom att kraftfullt och snabbt fördöma det faktum att Jörg Haiders främlingsfientliga och antieuropeiska parti deltar i den österrikiska regeringen , vilket saknar motstycke sedan andra världskrigets slut , har Europeiska unionen signerat sin politiska födelseakt och bekräftat att den inte endast är en ekonomisk och finansiell gemenskap , en stor marknad , " affärsmännens Europa " .
Just nu blottas en del av dess framtid , dess innersta väsen , dess själ .
För första gången har Europaparlamentet kunnat göra sin röst hörd .
De europeiska socialdemokraternas upprop , på Olivier Duhamels initiativ , har väckt sinnena och möjliggjort ett beslutsamt och direkt politiskt gensvar på denna helt nya och oacceptabla situation .
14 europeiska stater har gett prov på denna beslutsamhet genom att enhälligt och omedelbart - med A. Guterres röst - fördöma risken för en österrikisk politisk urspårning .
Detta modiga ställningstagande inleder ett nytt kapitel i det europeiska byggets historia .
Äntligen går vi tillbaka till ursprunget , en gemenskap uppbyggd på viljan att vända ryggen åt ett förflutet märkt av hat och utestängning och i stället ansluta oss till humanistiska värden som öppenhet och tolerans .
Europa hade förmågan att resa på sig och fördöma det oacceptabla .
Men med tanke på att det saknas juridiska instrument för denna politiska vilja - de sanktioner som föreskrivs i artikel 7 i fördraget är nästan omöjliga att tillämpa - kommer då Europa att kunna hålla huvudet högt inför hotet om en systematisk blockering av hela den institutionella strukturen ?
I dag gäller det Europas trovärdighet , innan vi i morgon kan ta emot de ännu sköra demokratierna i det f.d. östblocket .
Europa måste nu omsätta sina ord i handling för att i allas ögon bekräfta hur stora våra återfunna ambitioner faktiskt är . .
( FR ) När vi nu röstar om en gemensam resolution mot att nynazister skall ingå i en regering i Europeiska unionen , måste jag beklaga att kompromisstexten framför allt saknar bestämdhet .
Jag röstar för den , för det vore omöjligt att Europaparlamentet inte skulle ta ställning efter gårdagens mycket utmärkta politiska debatt .
Men personligen fortsätter jag att bekämpa extremhögern , jag fortsätter att samla in underskrifter till en petition för att kräva åtgärder som kan gå så långt som till att utesluta Österrike och jag fortsätter genom att organisera en stor medborgardemonstration i Lille på lördag kl .
15.00 .
Fascismen och nynazismen är som cancer !
Det djävulska djuret har väckts !
För mig är det inte tal om att låta dem utvecklas och frodas utan att slåss med stor energi .
Europa föddes ur en vilja till fred , frihet och tolerans .
Det kommer inte på fråga att Europa skall acceptera att hysa främlingsfientliga , rasistiska och antisemitiska ministrar .
Räkna inte med att jag förblir stum och passiv . .
( EN ) I gårdagens debatt i Europaparlamentet uttryckte en del parlamentsledamöter oro över att vi lägger oss i ett medlemslands interna angelägenheter .
En sådan oro är onödig .
Europaparlamentet har aldrig tvekat att kommentera en utveckling man inte samtycker till i medlemsstaterna .
Vi har fördömt baskisk och irländsk terrorism .
Vi har motsatt oss rasism och kränkningar av minoriteters rättigheter .
Det är vårt ansvar som parlament , särskilt som Europeiska unionens demokratiskt valda röst , att kritiskt kommentera den nuvarande politiska utvecklingen i Österrike , vilken står i konflikt med parlamentets linje .
Genom att kommentera och klargöra vår ståndpunkt hindrar vi inte något parti i Österrike att bilda en koalitionsregering .
Vi förklarar ändå för dem , vilket det är vår rättighet och plikt att göra , att ett sådant beslut , om de fortsätter på det sättet , kan leda till vissa konsekvenser och att vi i själva verket varnar dem på förhand .
Andra påstår att vi borde skjuta upp domen tills vi ser detaljerna av en sådan överenskommelse .
Ett sådant synsätt är inte bara en politisk smitning , det är uttryckligen farligt .
Genom att nå en överenskommelse med Jörg Haider och hans parti , skulle de österrikiska kristdemokraterna i ett slag ge högerextremismen politisk legitimitet och dessutom ge dem tillgång till makt - vilket de kommer att använda som startplatta för ännu större valframgångar .
Därför måste Europeiska unionen klargöra sin ståndpunkt beträffande den nuvarande situationen i Österrike . .
Vi har röstat för den gemensamma resolutionen för att uttrycka vår solidaritet med alla dem som utsätts för främlingsfientlighet och rasism .
Vi har också röstat för resolutionen i protest mot den avskyvärda politik Jörg Haider står för .
Vi är dock mycket kritiska till de metoder de 14 medlemsländerna använt sig av i denna fråga .
I resolutionen saknas en tydlig hänvisning till respekten för medlemsländernas nationella identitet och konstitutionella traditioner i enlighet med artikel 6 i fördraget .
Det saknas också en punkt om EU : s medansvar för den sociala och politiska utveckling i Europa och Österrike som varit en av förutsättningarna för Haiders valframgång .
Högerextremism är - idag , som tidigare i Europas historia - resultatet av otrygga sociala och ekonomiska livsvillkor .
Den nedskärningspolitik som följt i EMU-anpassningens spår har befrämjat högerextremismens framgångar .
En radikal politik för trygghet och rättvisa i varje land är den bästa garantin för en demokratisk utveckling i Europa .
Denna förklaring avger jag på CSU-gruppens vägnar .
Det är outhärdligt att EU blandar sig i regeringsbildningen i en medlemsstat .
Det tillkommer inte EU att göra så .
I stället för ett förhastat fördömande av FPÖ och den österrikiska regering som är under bildande fordras först och främst en kritisk undersökning och värdering av regeringsförklaringen och partiprogrammet samt koalitionens politik .
Först efter att med kritiska ögon ha satt sig in i den kommande politik som de i koalitionssamtal inbegripna partierna ämnar driva har man möjlighet att avgöra huruvida denna regering strider mot Europas demokratiska anda .
Detta betyder inte att vi sympatiserar med Haider .
CSU : s europeiska parlamentsledamöter hyser inga som helst sympatier för FPÖ-ledaren Haider .
Som politiker måste vi tvärtom ställa oss frågan varför 27 procent av den österrikiska befolkningen valde ett parti som FPÖ vid valen i oktober 1999 .
Vi måste analysera orsakerna till detta och försöka undanröja de orsaker som leder fram till sådana resultat .
Endast en analys av FPÖ : s argument och politiska innehåll kan förhindra en radikalisering av politiken i Österrike .
I Europaparlamentets resolution frågar man däremot inte efter orsakerna till det österrikiska valresultatet och pekar heller inte på några möjliga lösningar .
Detta är grunden till varför CSU : s Europagrupp uttalar sig mot resolutionen .
Det är med stor oro vi åser de tilltagande högerextrema krafterna i Europa , framför allt i Österrike , Tyskland , Frankrike , Belgien och Italien .
Det är mycket viktigt att diskutera dess djupare orsaker och att vidta nödvändiga åtgärder för att bekämpa dem .
Eftersom vi vet att ökade sociala klyftor , arbetslöshet , problem med fattigdom och social utslagning skapar misstroende bland medborgarna och skapar gynnsamma förutsättningar för den högerextrema populismen , är det mycket viktigt att de europeiska institutionerna vidtar nödvändiga åtgärder för att förhindra att de rasistiska och främlingsfientliga ideologierna går framåt .
Detta kräver djupa förändringar av den ekonomiskt sociala politiken i den nyliberala kapitalismen , en prioritering av åtgärder för att skapa kvalitetsanställningar med rättigheter , en politik för att stärka en demokrati där medborgarna deltar och en utbildning med särskild uppmärksamhet på demokratiska värden och solidaritet .
På samma sätt som vi fördömer och bekämpar högerextremismens idéer och verksamhet , uttrycker vi solidaritet med det österrikiska folket och vi stöder alla de krafter som för att fördjupa demokratin kämpar mot rasismen och främlingsfientligheten . .
( FR ) " Ty han visste det som den jublande skaran var okunnig om och som man kan läsa om i böcker , nämligen att pestens bacill aldrig vare sig dör eller försvinner , att den under decennier kan slumra i möbler och källare , koffertar , näsdukar och pappersluntor och att den dag måhända skulle komma , då pesten , människorna till olycka och varnagel , ånyo skulle väcka sina råttor och sända dem ut att dö i en lycklig stad . "
Med dessa ord avslutar Albert Camus en lång allegorisk berättelse som beskriver Oraninvånarnas svåra kamp mot pesten , för att efter andra världskrigets slut påminna oss om att kampen mot nazismen - " den bruna pesten " som den då kallades - inte kan krönas med en definitiv seger .
Att rashatet , det främlingsfientliga våldet , rädslan och avvisandet av det annorlunda alltid kan återuppstå och komma att dominera vilken grupp av människor som helst , eftersom det är något som bottnar i människans lägsta sidor .
Det är i denna bemärkelse de aktuella händelserna i Österrike måste betraktas som tragiska .
För första gången sedan andra världskriget står ett öppet pronazistiskt , rasistiskt och främlingsfientligt parti på tröskeln till makten i ett europeiskt land .
Inför detta hot - som i sig bär på ett förnekande av det europeiska byggets centrala idé - får ingenting stå i vägen : varken juridiska hårklyverier om vad fördraget tillåter och inte tillåter eller legitima frågetecken kring rätten till inblandning , eller en löjeväckande respekt för en formell demokrati , och framför allt inte den känsla av maktlöshet som griper oss inför en händelse som vi med våra övertygelsers fulla kraft vägrar att acceptera , men som vi inte har någon kontroll över .
Som förtroendevald från ett franskt utomeuropeiskt departement , La Réunion , en sammansmältningens och blandningens jordmån där befolkningen under de tre senaste seklerna har formats av successiva tillskott av européer , svarta från Afrika och Madagaskar , soldater från Indien och Pakistan och till och med kineser , upplever jag varje dag den djupaste sanningen i Saint-Exupérys ord : " Om du är olik mig , min bror , gör du mig inte illa , nej långt därifrån , du berikar mig ! " .
Det är den mänskliga mångfalden som har skapar vår främsta rikedom , och därför är det min plikt att förfölja och fördöma allt som kan kränka den - var den än visar sig .
Av alla dessa skäl har jag med stor beslutsamhet röstat för den resolution om den österrikiska regeringsbildningen som lagts fram i kammaren . .
( FR ) Jörg Haiders befordran , till följd av att FPÖ och den konservativa högern bildar regering , markerar en förfärande återuppståndelse av det monster som liberalismen skapat .
FPÖ : s framgångar har lika mycket att göra med de intyg om respektabilitet som tilldelats av den österrikiska högern och socialdemokratin som med de sistnämndas politik , vars sociala misslyckande har banat vägen för extremhögerns populism .
I resolutionen aviseras eventuella diplomatiska åtgärder för att politiskt isolera den nya regeringen , men här yppas inte ett ord om de bakomliggande orsakerna till fascismens uppgång .
Denna framgång kan förklaras av förvirringen bland de folk som fallit offer för penningdyrkan och av de ledande klassernas val att främja en kraftig åtstramning , för att hela tiden kunna driva svångrems- och avregleringspolitiken ett steg längre .
För att opponera oss mot det främlingsfientliga talet hos en diktatorlärling som längtar tillbaka till det tredje riket , är alla tillfällen bra för att uttrycka vår solidaritet med de antifascistiska österrikarna .
Därför kommer vi att rösta för denna resolution , trots de hycklande hänvisningarna till en " europeisk demokratisk modell " , som mer påminner om en fästning där man jagar , utvisar och låser in dem som lever under illegala förhållanden , när man inte sätter dit tonåringar . - ( DE ) Jag har just röstat mot resolutionsförslaget om Österrikes situation i betraktande av en möjlig regeringsbildning mellan Österrikiska folkpartiet ( ÖVP ) och Österrikiska liberala partiet ( FPÖ ) .
Jag håller det för kontraproduktivt att höja Jörg Haiders anseende som " Europas syndabock " - en allvarlig nynazist och ledande rasist .
Givetvis instämmer jag på intet sätt i denne högerpopulists publicerade uttalanden och fördömer på det starkaste all främlingsfientlighet och varje ansats till bagatellisering av Hitler-regimen .
Jag befarar dock att en blott och bart emotionellt präglad reaktion från Europa på vad som sker i Österrike kommer att mångfaldiga Haiders anhängare .
Europeiska unionen får inte skänka honom en PR-effekt som annars inte kan fås för pengar .
FPÖ : s styrka kan härledas till svagheten hos dem som hittills har regerat .
Här bär de österrikiska socialisterna huvudansvaret .
Först efter att utan framgång ha propagerat hos FPÖ för accepterandet av en minoritetsregering och uppenbarligen förgäves ha erbjudit FPÖ ministerposter påbörjade Österrikiska socialdemokratiska partiet ( SPÖ ) sin massivt förda kampanj mot Haider .
Den hotande maktförlusten döpte de om till en " heroisk kamp för upprätthållandet av värderingar " och helt enkelt ett omedelbart förestående " avgörande mellan demokratins vara eller icke vara " .
Detta är en smädelse mot väljarna i mitt grannland , vilken jag inte kan ställa upp på .
Vi tyska kristdemokrater valde en annan strategi i kampen mot extremister och tog i klartext avstånd från dem .
Vi avslöjade de innehållsliga bristerna hos REP ( " die Republikaner " ) , vilka visade sig vara nationalistiska , främlings- och minoritetsfientliga .
I dag saknar REP representation i de flesta kommunalparlament .
Den tyska vägen är ingen garanti för att denna radikala rörelse inte växer sig stark på nytt .
Den kan inte tillämpas var som helst , eftersom varje medlemsstat har sina egna villkor .
ÖVP ( Österrikiska folkpartiet ) , som man inte längre kan ignorera ens på europeisk nivå , vågar sig på försöket med en koalition , för det österrikiska styrets skull .
Detta kan lyckas endast om man träffar överenskommelser som på ett övertygande sätt bottnar i viljan att upprätthålla demokratiska grundläggande värderingar .
Rådet har blandat sig i oöverlagt , utan att invänta resultaten av koalitionsförhandlingarna eller ett regeringsprogram .
Detta fördömande är precis lika litet acceptabelt som hotet om att bryta kontakterna med republiken Österrike En väl befäst demokrati kräver att man är vaksam och inte blundar med ena ögat .
Vi måste reagera offensivt och med argument mot radikala personer såväl från höger som från vänster .
Jag skulle ha önskat mig samma häftiga europeiska protest när socialisterna såg sig redo att göra gemensam sak med efterföljarna till den människoföraktande och människoförföljande regimen i DDR .
Sedan dess bildar de regering i olika tyska förbundsländer .
Jag instämmer helt och fullt i de redogörelser som Europeiska kommissionens ordförande Prodi lämnade under dagens sammanträde .
Han talade om vår plikt att inte isolera medlemsstater utan att göra allt för att knyta dem till gemensamma europeiska värderingar . .
( FR ) Jag har röstat emot den gemensamma resolutionen om situationen i Österrike .
Österrike är en fri , oberoende och suverän nation .
Följaktligen kan varken rådet , kommissionen eller Europaparlamentet blanda sig i en medlemsstats interna organisation .
Valen i Österrike har genomförts på ett fritt , regelmässigt och demokratiskt sätt .
Därför är EU-institutionernas inblandning i det här landet oacceptabelt ; det är en kränkning av det europeiska fördraget ( artikel 7 i Amsterdamfördraget ) .
Likväl har dessa institutioner inte tvekat om att godkänna Turkiets anslutning till Europeiska unionen , samtidigt som man känner till att det förekommer kränkningar av de mänskliga rättigheterna .
Ingen händelse av ett sådant slag har inträffat i Österrike .
Detta prejudikat , som skapats på initiativ av det portugisiska ordförandeskapet , är oroväckande för Europeiska unionens framtid : dels avslöjar den politiska bannlysningen av Österrike att likriktningen har ett oroande övertag , och dels kommer själva demokratins princip att förstöras om regeringarna i Europeiska unionens medlemsstater i framtiden först måste - inte få folkets förtroende - utan nomineras av överstatliga organ .
Kommer det att ens vara lönt att anordna val under sådana omständigheter ?
Det är inte så man skapar förutsättningarna för att Europas nationer skall kunna leva i harmoni och samarbeta för en gemensam framtid .
Jag röstar emot det gemensamma resolutionsförslaget angående resultatet av valet i Österrike och förslaget att bilda en koalitionsregering mellan ÖVP och FPÖ av tre olika skäl : för det första därför att man inte gick med på varken de separata omröstningar vi krävde eller några av de föreslagna ändringsförslagen , vilka i sin helhet skulle ge texten en annan samstämmighet och mening ; för det andra för att den resolution som nu godkänts innehåller en motsägelse i själva texten : å ena sidan , i skäl D erkänner man att EU : s och dess institutioners betoning av främjandet av försvaret av de europeiska demokratiska värdena innehåller ett erkännande av Österrikes folks och den österrikiska statens demokratiska rättigheter och konstitutionella privilegier , och å andra sidan , tillåter man sig , och till och med gratulerar ( punkt 4 ) till de politiska avsikterna med det portugisiska ordförandeskapets uttalande , vilket inte , enligt vår mening , var mer än en förhastad , olycklig och obefogad inblandning i Österrikes folks och den österrikiska statens demokratiska rättigheter och konstitutionella privilegier ; vi förstår det så , och detta är det tredje skälet till vår röst , att resultatet av Österrikes fria och demokratiska utövande av rösträtten inte kan dömas , det skall respekteras eller åtminstone skall man inte döma det på förhand , vilket sker i detta fall .
Faktum är att med denna resolution och övriga liknande ståndpunkter , visas inte minsta hänsyn till den uttalade viljan hos väljarna i en av EU : s medlemsstater , förutom att EU inte tolererar ( lustigt nog i toleransens namn ) att regeringslösningen som detta resultat gav upphov till går sin egen väg och får bevisa sina upprepade avsikter och politiska förslag främst inför de anklagelser den utsätts för .
Resolutionen gör också att man på ett dumt sätt genom manipulation och genom att göra dem man vill fördöma till offer , stärker deras ställning och till slut får ett mycket allvarligt precedensfall , inom själva EU .
Detta kan bara leda till ett växande undergrävande av det förtroendefulla klimat och den ömsesidiga respekt som bör råda mellan nationer och medborgare vilka i en anda av likhet och respekt för den nationella suveräniteten vill fortsätta på en gemensam väg .
Den väg på vilken de liksom vi står i motsatsställning till rasistiska och främlingsfientliga ståndpunkter som grasserar litet överallt i Europa , men som föredrar att på ett beslutsamt sätt angripa de orsaker som har gett upphov till dem . .
( FR ) Den omröstning som just har ägt rum här är historisk , för det är första gången som vi med en så stor oro diskuterar den interna politiska situationen i en av våra medlemsstater .
Jag tror det är lämpligt att frågan om institutionella principer och regler ställs åt sidan .
Jag uppmuntrar rådet och dess ordförandeskap att fortsätta försvara unionens grundläggande värderingar .
Och jag uppmanar kommissionen att vara mindre försiktig .
Med denna resolution tar parlamentet sitt ansvar .
Men samtidigt är den resolution som i dag antagits i mina ögon ett minimum minimorum , det minsta vi kan göra .
Personligen har jag försvarat en ännu hårdare ståndpunkt och därmed stött ändringsförslagen 1 , 4 , 6 , 7 , och 8 , såväl som det muntliga ändringsförslag vilket föreslogs av socialistgruppen .
Jag tror faktiskt att det är en nödvändighet att rådet endast accepterar tekniska förbindelser med företrädare för den österrikiska regeringen , där FPÖ-medlemmar kommer att ingå .
Att låta Jörg Haiders parti ingå i en regeringskoalition kommer att banalisera extremhögern i Europa , och utgör ett ytterst allvarligt prejudikat som skulle kunna dra med sig andra unionsmedlemmar eller kandidatländer .
Här tar det österrikiska konservativa partiet ett historiskt ansvar .
Det är våra grundläggande värden som står på spel ; i egenskap av européernas demokratiskt valda företrädare har vi inget val .
Vi måste , våra väljare kräver det , vägra det oacceptabla .
När barbariets spöke dyker upp igen skall vi veta följande : " Att inte opponera sig är att kapitulera " . .
( FI ) Jag röstade blankt vid omröstningen om resolutionen .
Jag fördömer Jörg Haiders rasistiska och främlingsfientliga linje .
Jag kan emellertid inte acceptera att EU : s organ gör en politisk intervention i en medlemsstats inrikespolitik .
Därför kan jag varken godkänna punkt 4 i den gemensamma resolutionen eller rösta för resolutionen , inte ens mot extremhögern . .
Det är uppenbart att de politiska ledarna i Europa har rätt och skyldighet att reagera mot Haider och hans parti .
De politiska ledarna i Europa har rätt att uttala sin uppfattning om den politiska utvecklingen i ett annat medlemsland , på samma sätt som en statsminister kan uttala sig om rasistiska politiker i en kommun .
Den finländska erfarenheten är emellertid att integrering är ett bättre sätt att bekämpa antidemokratiska krafter än att isolera .
Därför röstade jag emot punkt 2 i resolutionen .
Detta förutsätter dock att alla parter respekterar mänskliga rättigheter .
EU-ordförandeskapets " gemensamma reaktion " på regeringsbildningen i Österrike är juridiskt felaktig .
De 14 medlemsländernas reaktion saknar stöd i fördragen .
Vi skall inte heller isolera de krafter i Österrike som vill arbeta för mänskliga rättigheter .
Trots dessa mina invändningar mot rådets agerande och min åsikt att det är bättre att verka för integrering än genom isolering , var det viktigt att visa klart var Europaparlamentet står i frågor om rasism , varför jag röstade för resolutionen i slutomröstningen .
Härmed avslutas omröstningarna .
 
Avbrytande av sessionen Jag förklarar Europaparlamentets session avbruten .
( Sammanträdet avslutades kl .
12.25 . )
