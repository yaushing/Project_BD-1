 
Justering av protokollen från de två föregående sammanträdena Protokollen från sammanträdena torsdagen den 3 februari och måndagen den 14 februari har delats ut .
Protokollet från den 3 februari delades i själva verket ut redan i Bryssel .
Det är kanske därför som en del kolleger inte hade fått det .
Finns det några synpunkter ?
( Prokollet justerades . )
Fru talman !
Jag brukar alltid vara här när sammanträdet inleds på måndagarna klockan 17.00 .
I går var det dock omöjligt för mig och för många andra europeiska ledamöter att närvara , eftersom Air France-flyget som brukar ta oss hit , 14.15-flyget , ställdes in utan några förklaringar från flygbolagets sida , och därför var klockan mycket när vi kom fram .
Om Air France fortsätter att bojkotta Europaparlamentet , bör åtgärder vidtas för att förhindra en upprepning av detta .
( Applåder ) Tack , herr Medina Ortega .
Jag delar fullt ut det beklagande som ni uttrycker .
Skulle ni vänligen vilja skriva till mig så att jag med stöd av bevis kan anmäla detta till de behöriga ansvariga såväl hos Air France som den franska regeringen ?
Jag tror verkligen att det inte längre är möjligt och att vi absolut måste protestera med full energi .
Fru talman !
Igår upplevde jag och Medina Ortega samma sak .
Jag tycker att de franska myndigheterna - som har äran att hysa Europaparlamentets säte i Strasbourg - bör vara medvetna om sitt ansvar för att garantera fungerande kommunikationer med alla unionens huvudstäder .
Just det , herr Napolitano , tack för det .
Fru talman !
Det handlar här inte om försenade plan : jag skulle vilja be om ursäkt för min kollega i Gruppen De gröna , Caroline Lucas , som är brittisk ledamot .
Hon kunde inte närvara eftersom hon hade arresterats vid en demonstration mot kärnkraft i Glasgow i går morse .
Hennes identitet noterades : det framkom mycket tydligt att hon är ledamot av Europaparlamentet , ändå kvarhölls hon i arrest hela dagen .
Jag anser att det är absolut oacceptabelt och jag ber er - jag har för övrigt skrivit till er tillsammans med min kollega Hautala i det avseendet - intervenera hos de brittiska myndigheterna för att sådana händelser inte skall upprepas och att man ber Lucas om ursäkt .
Tack , herr Lannoye .
Jag har fått er skrivelse och har redan vänt mig till den brittiska delegationen .
Fru talman !
Med tanke på omröstningen i dag vill jag be om något som jag berörde redan i går vid debatten om Equal-betänkandet .
Jag ber om att man uppskjuter omröstningen i dag om gemenskapsinitiativet Equal , eftersom vi helt enkelt behöver litet mer tid för att komma överens om en viktig punkt .
Jag är optimistisk och ser verkligen med lugn och tillförsikt fram emot omröstningen ; vi kommer att få ett synnerligen brett godkännande av detta yttrande om Equal .
Vi behöver bara litet mer tid för att utarbeta detaljerna i samband med asylfrågan , och jag ber därför om att omröstningen genomförs i morgon i stället för i dag .
Fru talman !
För att fortsätta från den punkt som Lannoye tog upp : Lucas arresterades precis utanför Glasgow för att hon protesterade mot Tridentbasen i Faslane .
Jag sympatiserar mycket med den protesten .
Jag har dock ingen sympati för Lucas som försöker gömma sig bakom sin parlamentariska immunitet .
Jag har också varit arresterad för att ha protesterat i Faslane .
Jag gömde mig inte bakom någon immunitet .
Jag tog det straff som jag fick .
Lucas borde göra detsamma .
Fru talman !
Jag skulle vilja kommentera Stenzels yrkande om att skjuta upp omröstningen om gemenskapsinitiativet Equal till i morgon .
Detta initiativ har faktiskt diskuterats mycket livligt i utskottet , och eftersom det är ett viktigt förslag från kommissionen , som gäller de överenskommelser vi träffade förra året , tycker jag att det kan antas .
Vi är överens med Stenzel om att yrkandet om uppskjutande kan bifallas för att finna största möjliga samförstånd mellan grupperna , så att parlamentet med bredast möjliga majoritet uttrycker sin ståndpunkt om detta initiativ .
Finns det några kolleger som vill yttra sig mot Stenzels begäran , som Ghilardotti just stödde ?
Eftersom det inte är så , tar vi upp den till omröstning .
( Parlamentet gav sitt samtycke . )
Fru talman !
Enligt artikel 29.4 skall ni hållas informerad av de politiska grupperna om varje ledamot som anslutit sig till en ny politisk grupp eller lämnat en politisk grupp .
Har ni fått någon anmälan om att några medlemmar lämnat gruppen Europeiska folkpartiet eller tillhör Österrikiska folkpartiet fortfarande denna politiska grupp ?
Herr Corbett , jag har inte hört talas om någonting .
Fru talman !
Jag är mycket förvånad över denna reaktion från kollegan Corbett .
Han borde söka andra möjligheter för att profilera sig , än att här yttra sig om en sådan punkt !
( Applåder ) Vi är solidariska med våra österrikiska vänner , som tidigare har visat sig vara goda européer .
Ni har vårt fulla stöd !
( Applåder )
 
Föredragningslista När det gäller föredragningslistan för torsdagen föreslår jag er , mot bakgrund av en begäran som inlämnades i går vid plenarsammanträdet , att förlänga debatten om brådskande och aktuella frågor med en halvtimme , det vill säga fortsätta fram till kl .
18.00 .
Omröstningen kommer att äga rum kl .
18.00 .
( Parlamentet gav sitt samtycke . )
 
Strategiska mål och lagstiftningsprogram från kommissionen Nästa punkt på föredragningslistan är den gemensamma diskussionen om kommissionens uttalanden om sina strategiska mål för en femårsperiod och om det årliga lagstiftningsprogram för år 2000 .
Jag ger genast ordet till ordförande Prodi .
Fru talman , ledamöter !
Ett femårsprogram är ett viktigt åtagande och därför tyckte jag det var bättre att ni alla fick hela texten till talet utdelad , den finns på fyra språk .
För att respektera tidsbegränsningen skall jag endast ta upp de stora dragen i mitt program : ett program för början av en mandatperiod och för början av ett nytt sekel under vilket man har både rättighet och skyldighet att se Europa i ett vidare perspektiv , ett Europa som för närvarande upplever en motsägelsefull tid .
Vi skall komma ihåg att Europa under sina femtio års historia har gett oss fred , säkerhet och frihet , och att det enade Europa också har bidragit till att ge oss en period med aldrig tidigare skådat välstånd .
Nu känner vi av början på en solid återhämtning som även verkar kunna bli mycket varaktig om vi för en klok politik , en återhämtning som är en logisk följd av de ansträngningar vi har gjort .
Vi får den inte gratis , utan som en konsekvens av saneringen av de offentliga finanserna i Europas länder , som har hållit inflationen under kontroll med en klok politik inriktad på kostnadskontroll och ökad produktivitet .
Detta i ett Europa som har inlett en energisk omstrukturering av sina industrier , banker och sin offentliga service , även om denna process ännu inte är fullbordad , även om det fortfarande är långt kvar att gå .
Trots dessa aspekter finns det ändå besvikelse och oro i Europa : besvikelse och oro för arbetslösheten som inte minskar tillräckligt snabbt , för en teknisk eftersläpning som framstår som större och större , och som framför allt börjar åtföljas av en kraftig eftersläpning också inom det vetenskapliga området , för de europeiska institutionerna som verkar vara långt efter , som inte verkar vara tiden vuxna , i första ledet kommissionen själv .
Kommissionen kris var faktiskt en avgörande punkt i förhållandet mellan Europa och dess medborgare , och det låga valdeltagandet i Europavalen var ett oroande tecken på detta .
Något som går ännu djupare är dock känslan av osäkerhet , känslan av att inte vara förberedd för den nya värld som växer fram , en värld som förändras totalt , som genom globaliseringen kommer att förändra också våra referensramar .
Detta är ingenting alldeles nytt i historien : Europa har redan tidigare en gång genomgått en liknande förändring med en explosionsartad ökning av marknaderna , förändrade referensramar och en ny världsuppfattning .
Jag syftar på femtonhundratalet , efter upptäckten av Amerika , då allting förändrades .
Vissa länder - såsom Frankrike och Spanien - visste att svara på utmaningen och gav upphov till stora nationalstater .
Andra länder - såsom Italien - klarade inte denna utmaning och förlorade all den dominans de hade byggt upp under millenniets första hälft : en dominans inom vetenskap , teknologi , ekonomisk utveckling , försvarsstrukturer och militär organisation , filosofi och litteratur .
I dag står Europa inför en liknande utmaning och vi vet att historien kommer att vara lika skoningslös som förr i tiden .
Mot bakgrund av dessa stora förändringar fordras ett ekonomiskt starkt Europa för att förhindra att våra nationalstater även nu försvinner genom en globalisering med dimensioner och utmaningar utan motstycke i vår historia .
Globaliseringen påbjuder nämligen enhet .
Varje dag hör vi nyheter om nya avtal på global nivå och varje dag hör vi nyheter om förändringar också på europeisk nivå .
Men ännu mer nödvändigt är att Europa känner sig starkt på det politiska planet .
Tidigare har den inre marknaden och den gemensamma valutan varit den fasta punkten i vårt handlande , det bärande elementet i Europas liv .
I dag är de nya gränserna för den europeiska integrationen politiska gränser : den gemensamma utrikes- och säkerhetspolitiken , den inre rättvisan och säkerheten och - på ett underordnat plan - den avgörande frågan om de grundläggande politiska värderingar vår samexistens vilar på .
Därför har kommissionen antagit den strategiska planen för 2000-2005 , en plan som genast översändes till Europaparlamentet , som ni redan känner till och som jag alltså inte skall beskriva i detalj här .
Någon kanske anser att den är för allmänt hållen , men inga politiska instanser upprättar detaljerade femårsplaner .
Detta är Europeiska unionen , inte Sovjetunionen .
I vår plan anges de stora referensramarna , vår verksamhets inriktning i stort : för det första att utveckla nya styrelseformer för Europa , för det andra att expandera och utvidga området för fred , frihet och säkerhet , för det tredje att lansera en ny ekonomisk utvecklingsfas , för det tredje att värna och öka livskvaliteten .
Dessa är våra stora handlingslinjer för de kommande fem åren .
Vad den första beträffar - de nya styrelseformerna för Europa - vet ni redan att kommissionen har åtagit sig att lägga fram en vitbok och inte en komplett lagtext eftersom kommissionen inför de stora frågor som förändrar strukturen för vårt umgänge först tar fram ett debattunderlag .
Sedan diskuterar vi innehållet med er , och ur detta uppstår ett först politiskt dokument och slutligen en lagtext .
Detta är ett öppet och kraftfullt sätt att gå till väga , så att alla europeiska institutioner och Europas befolkning involveras .
Denna vitbok är ett svar på de utmaningar utvidgningen ställer upp .
Det är utvidgningen som tvingar oss att se över hur alla våra institutioner fungerar , att till och med se över vår politik - all vår politik - och framför allt tänka igenom vad vi skall fortsätta att göra på unionsnivå när medlemsländerna är tjugofem eller trettio , vad som bättre görs av de enskilda staterna , regionerna eller de lokala myndigheterna .
Men det är inte bara utvidgningen som driver oss till denna översyn : som jag sade nyss är det också globaliseringen av ekonomin och politiken .
Vi måste styra Europa så att vi blir mer effektiva , kommer närmare medborgarna och verkar för allas delaktighet .
Först och främst måste vi ta itu med den stora frågan om kvinnors delaktighet .
I den jämförelse mellan Europa och Förenta staterna som nyligen gjordes är en av de stora skillnaderna inte så mycket arbetskraftens rörlighet eller tillgången på riskkapital utan kvinnors deltagande i det ekonomiska livet , ett deltagande som i Förenta staterna har helt andra dimensioner än i Europa .
Det handlar om ett område där Europa tvärtom alltid har varit ledande : detta måste vi alltså tänka igenom på djupet och öppet , och alla institutionerna - kommissionen , parlamentet och rådet - måste tänka igenom sin roll och sin politik .
Vi kommer alltså att omedelbart börja arbeta med denna vitbok , även om vi måste avvakta resultaten fån regeringskonferensen innan vi slutför den och den därför inte kan läggas fram förrän våren 2001 .
Det blir ingen filosofibok utan en konkret bok med många detaljerade förslag .
Vi - kommissionen - är de första att veta att vi måste göra en total översyn av oss själva , och därför kommer vi att göra två saker : vi kommer att engagera oss och vi engagerar oss redan nu till fullo i den interna reformen , och vi kommer att tänka igenom vår politik på djupet .
Jag har bett alla kommissionärer - och vi kommer att be dem om en ännu djupare analys - att identifiera all verksamhet som kan läggas ned .
Kommissionen måste fastställa sin kärnverksamhet , den verksamhet vi skall koncentrera oss på , och upphöra med mindre viktig verksamhet för att frigöra nya resurser och få ett korrektare och mer samarbetsbetonat förhållande med de enskilda länderna , med regionerna och med de lokala samhällena .
Vi skall alltså frigöra nya resurser , men det kommer också en tid - fruktar jag , och jag vill säga det här inför parlamentet - då även dessa nya resurser som vi redan håller på att frigöra inte kommer att vara tillräckliga för att vi skall kunna ta itu med våra nya uppgifter : jag tänker på utvidgningen , på den nya rättsliga och inrikespolitiska sektorn , på hälso- och sjukvårdsfrågorna , på miljöfrågorna .
Den dagen , när vi har utnyttjat alla våra resurser maximalt , kommer jag inte att tveka att inställa mig inför er för att be om nya resurser , men jag säger redan nu att om vi inte har erforderliga resurser måste vi vägra ta på oss några nya uppgifter , eftersom det inte finns någon överensstämmelse mellan de nya uppgifter vi tar på oss och de resurser vi har till vårt förfogande .
Vad den interna reformen beträffar känner ni väl till det engagemang min kommission har lagt ned på denna fråga från första dagen .
Jag vet mycket väl att vi inte kan uppnå några politiska mål om kommissionen inte reformerar sig internt kraftigt och genomgripande , om vi inte blir effektivare , om vi inte tar ett effektivitetssprång inom alla sektorer med början i den sektor där vi hittills har samlat på oss den mest dramatiska eftersläpningen , det vill säga inom det externa biståndet .
Att ge hjälp snabbt när den behövs räddar människoliv .
Att ge den för sent kan i många fall vara värre än att inte ge den alls .
När jag talar om externt bistånd går mina tankar i första hand till Balkan , där det finns en stråle av hopp tack vare våra funktionärers engagemang på fältet , ett extraordinärt engagemang med tanke på de organisatoriska problem vi har .
Jag tänker även på Bernard Kouchners bemödanden , på stabilitetspakten som vi står bakom med kraft , med total hängivelse , men jag tänker också på de nya händelserna i till exempel Kroatien , där situationen har förändrats på några veckor : de europeiska institutionerna öppnade omedelbart dörren för en dialog med detta land , de mottog denna nyhet väl medvetna om att inte bara Bosniens utan framför allt Serbiens problem endast kommer att kunna lösas om vi slår en demokratisk järnring kring Serbien .
Detta är det nya element vi måste bidra till att införa på Balkan .
Vi måste bli effektivare på detta område , vi måste öppna Donau för trafik igen .
Det är motsägelsefullt att erbjuda hjälp till Rumänien och Bulgarien och låta dessa länders stora resurs vara blockerad .
Vi måste rena floden och därför kommer den miljöansvariga kommissionären under de närmaste dagarna att lägga fram detaljerade projekt för att få bukt med detta allvarliga problem .
Vi har gjort mycket på Balkan : den nya Europeiska byrån för återuppbyggnad av Kosovo , insatsstyrkan för Balkan , en ny förordning för att snabba upp rutinerna .
Vi måste dock absolut göra mer .
Vi måste liberalisera handelsutbytet inom regionen och utbytet mellan denna region och Europeiska unionen .
Vi måste bidra till att konstruera infrastruktur som bryter en sekellång isolering .
Vi måste intensifiera ansträngningarna för att i dessa länder bygga upp demokratiska och pluralistiska samhällen med ett civiliserat samhälles institutioner , offentliga strukturer , ordningsmakt och organisation , men framför allt måste vi få dessa länder att arbeta tillsammans och se regionen som en enhet både politiskt och ekonomiskt .
Om vi inte gör det har vi misslyckats med vår uppgift .
Minns att Marshallplanen på sin tid inte bara hade effekt på grund av sina stora resurser : den fick ännu större effekt eftersom den tvingade oss européer att arbeta tillsammans med ett nytt perspektiv , att ge vår politik och vår ekonomi en ny horisont .
Detta är vad vi måste göra för Balkan .
Europa måste för Balkanländerna och hela resten av världen bevisa sin förmåga att utvidga området för säkerhet , fred och frihet , sin kapacitet att spela en huvudroll på den internationella scenen .
Självfallet kommer vi åter igen tillbaka till utvidgningen , som måste genomföras genom att man samtidigt utvidgar området för säkerhet , fred och frihet .
Vi har lovat mycket i denna riktning men jag tror att vi kommer att kunna hålla våra löften även om vi har en mycket delikat uppgift framför oss .
Utvidgningen , som kommer att följa oss under hela vår femårsperiod och även senare - jag tänker på kandidatländernas förhoppningar - måste komma till stånd med säkerhet och objektiva kriterier , men den måste också komma till stånd så att man lugnar den allmänna opinionen i de berörda länderna och , än mer , lugnar vår egen allmänna opinion .
Det kommer att bli vänskap , harmoni och öppenhet , men också stränghet i utvidgningen .
Jag upprepar : vi måste lugna den allmänna opinionen i de länder som vill bli medlemmar , men vi måste lugna vår egen allmänna opinion ännu mer .
Våra skyldigheter upphör inte med utvidgningen , de upphör inte med Balkan .
Det finns några andra frågor som är avgörande : förhållandet med Ukraina , förhållandet med Ryssland , förhållandet med våra grannländer och i än högre grad den stora frågan om förhållandet med södra Medelhavsområdet , som kommer att bli den avgörande punkten i den europeiska historien , för kommande generationers säkerhet och trygghet i Europa .
I denna mening har vi en skyldighet mot hela Afrika : Afrika som man har vänt sig till med förhoppningar på den senaste tiden , som har fått mottaga erbjudanden men där ännu ingenting konkret har genomförts .
Afrika där övergången under de senaste åren inte har varit från totalitära regimer till demokrati utan tvärtom , från demokrati till totalitära regimer .
Afrika som är bekymmersamt för oss att konfronteras med .
Därför har vi ytterligare en uppgift på det internationella planet , vilken kommissionären med ansvar för handelsfrågor redan har föreslagit : uppgiften att återuppta Millennium Round , med ett stort tillmötesgående som vi redan tagit på oss och erbjöd redan innan Seattle , men som inte kunde konkretiseras .
Att alltså ta över bördan för vissa grundläggande problem från de fattigaste länderna , inte bara vad gäller avskrivning av skulder utan även att ensidigt öppna för handel med världens fattigaste länder .
Det krävs en ny lösning , annars kommer händelser som de i Seattle alltid att upprepas och förhindra att Europa utövar en positiv roll i historien .
Överallt i världen måste Europas agerande styras av stor respekt för principerna om frihet , respekt för individens rättigheter och respekt för minoriteters rättigheter .
Låt oss komma ihåg att vi , Europeiska unionen , är en union av minoriteter : alla vi är i minoritet i Europa .
Det finns en oro även hos våra femton länder , en oro som kanske kommer att uppstå igen under den kommande tioårsperioden .
Jag talar om fallet Österrike , där kommissionen har varit sin roll trogen .
Vi har verkat för sammanhållning av unionen men varit orubbliga i vårt försvar av fördragen , redo att bestraffa varenda litet övertramp som innebär ett brott mot principerna om demokrati , rättigheter och respekt för minoriteter .
Vissa har kritiserat mig för det lyckönskningsmeddelande jag skickade till kansler Schüssel .
Jag skall säga er : förväxla inte en nödvändig och pliktskyldig formell hövlighet med mindre reell fasthet .
Läs brevet igen : hänvisningen till unionens grundläggande värderingar är ett utdrag ur fördragets artikel 6 , jag upprepar artikel 6 i fördraget , och detta är ingen tillfällighet .
Jag frågar er också : tror ni att kommissionen någonsin har påmint någon annan nyvald europeisk regeringschef om dessa principer ?
Det är detta vi vill göra : bibehålla vår roll av övernationell struktur , bibehålla den roll vi har fått genom fördragen , men också vara obevekliga om principerna och utgå från fakta i våra bedömningar .
I november förra året lade kommissionen fram ett förslag till direktiv mot rasismen .
Jag ber rådet att snabbt anta det och jag ber parlamentet att hjälpa oss i denna kamp , som ytterligare fördjupar den grundläggande basen för vår sociala sammanhållning .
Jag skall avsluta med att snabbt påminna om de sista två punkterna i vårt program : ekonomin och livskvaliteten .
Jag har redan talat om ekonomin : vi är väl medvetna om vilka grundingredienserna är för att föra in Europa på vägen mot en återhämtning som kan vara länge och äntligen skapa arbetstillfällen .
Vi måste fortfarande hålla inflationen nere , fortsätta med avregleringen , värna konkurrensen i än högre grad , driva på spridningen av informationsteknologi och av all ny teknik , driva på vetenskapen , vetenskapens förfront , njuta av att befinna oss i vetenskapens förfront .
Det kommande toppmötet i Lissabon om dessa frågor - spridning av teknik och sysselsättningen - blir ett avgörande toppmöte .
Det behövdes fyra år innan vi kunde ha ett toppmöte av detta slag .
Nu kommer vi äntligen att ha det : vi får inte missa tillfället .
Det sista åtagandet är slutligen att öka livskvaliteten .
Vi inledde detta kapitel med vitboken om livsmedelssäkerhet : nu måste vi göra stora framsteg på miljöområdet .
Fallet med fartyget Erika och giftutsläppet i Donau visar hur angeläget det är med insatser på europeisk nivå till skydd för miljön .
Det är dags att fundera på , och sedan förverkliga , en europeisk räddningstjänst .
I allt för många fall hör man krav på detta efter det att katastrofen har inträffat .
Jag tror att man måste börja tänka på dessa saker innan katastroferna inträffar .
Dessa är de utmaningar vi har framför oss : vi som kommission men också alla de andra europeiska institutionerna .
Ledamöter , fru talman , hur skall vi mäta våra fem verksamhetsår ?
Hur skall vi mäta resultaten av dessa fem år ?
Jag vet inte , men en måttenhet kan helt klart vara den kamp vi måste utkämpa tillsammans .
Låt oss ta en mycket enkel parameter : valdeltagandet vid nästa Europaval .
Om det blir högre än vid det föregående valet betyder det att vi har vunnit vår kamp .
Fru talman , ärade ledamöter !
Vi har alla dessa stora politiska utmaningar framför oss , men vi har också stora möjligheter framför oss , just på grund av den återhämtning som har inletts .
Detta , ärade ledamöter , kan bli Europas decennium .
Jag säger : detta måste bli Europas decennium .
Fru talman , herr kommissionsordförande , kolleger !
Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater välkomnar denna debatt , och vi är positiva till att kommissionen har lagt fram ett dokument för att förbereda debatten .
Vi välkomnar också de slutsatser som vi finner i detta dokument .
Vi är i stora drag även positiva till talet som kommissionsordföranden Prodi just har hållit .
I slutsatserna i dokumentet står det att Prodi-kommissionens femåriga mandattid kommer att bli en tid av stora förändringar .
Europas integration kommer att fortsätta , och samtidigt kommer unionen att inleda en utvidgningsfas , som slutligen kommer att leda till en återförening av vår kontinent .
Det är anspråksfullt , ambitiöst , man kunde rent av säga att det är profetiskt .
Vi önskar er , herr kommissionsordförande , att detta kommer att lyckas .
Men vi säger också att nutiden är grundvalen för framtiden , och framtiden kommer vi bara att kunna gestalta om vi kan hävda oss i nutiden .
Det säger jag på allvar , och jag säger det med oro !
Med detta kommer jag in på den aktuella diskussionen beträffande de konflikter som för närvarande finns i Europeiska unionen .
Vi är en gemenskap inom Europeiska unionen .
Vi hör ihop , även om vi har problem .
Nu är det inte dags att isolera sig utan att knyta samman och gemensamt slutföra detta arbete med att ena Europa !
( Applåder ) Herr kommissionsordförande , ni har under de senaste veckorna alltid företrätt och försvarat Europaparlamentet .
Ni har uppfattar er som fördragens väktare - vilket är er roll .
Vi vill därför uttryckligen visa er vår respekt , vårt erkännande och vårt stöd , också för den av er nämnda skrivelsen till Republiken Österrikes förbundskansler .
( Applåder ) Herr kommissionsordförande , vi är ense med er när det gäller målsättningen : Vi vill ha ett starkt , handlingskraftigt och demokratiskt Europa under 2000-talet .
Ett Europa som försvarar sina värderingar beträffande den mänskliga värdigheten , demokratin och rättsstaten både inåt och utåt , och samtidigt iakttar sina intressen i världen med värdighet , tålamod och övertygande självmedvetande .
Europas , Europeiska unionens budskap till världen får inte vara förmätet eller rentav europeiskt nationalistiskt , nej , det måste innebära samarbete , partnerskap och fredlig utveckling .
Därför betyder globalisering för oss en chans att utforma denna enda värld , som krymper allt mer samman , i fredlig konkurrens och i solidaritet .
Sett på så vis innebär globalisering mer chans än risk , den för samman snarare än den skiljer åt , den innebär mer ömsesidigt berikande än avgränsning .
Men vi vet också att vi bara som européer , gemensamt , kan utforma dessa stora utmaningar i samband med globaliseringen .
Globalisering är inte bara en ekonomisk utan också en kulturell process .
Därför säger vi att vi vill ha partnerskap i världen , vi vill inte - som många förutspår - ha en kollision mellan kulturerna , en clash of civilisation , utan vi vill ha partnerskap , möten , utbyte och fred .
Men vi säger också att vi vill försvara detta europeiska samhälle av tolerans , och därför är en gemensam utrikes- , säkerhets- och försvarspolitik så viktig .
I dag börjar förhandlingarna med sex stater i Centraleuropa .
Därigenom sluter sig den europeiska familjen litet närmare samman .
Vi anser att det är riktigt , det som ni sade om Barcelona-processen : Alla länder i Medelhavsområdet måste erkänna den mänskliga värdigheten , demokratin och rättsstatligheten .
För oss , Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater , är det under de närmaste fem åren inte bara betydelsefullt med reformen av Europeiska unionens institutioner , utan också att vi bekänner oss till en gemensam valuta , och stabilitetspolitiken måste vara grundvalen för en konsolidering av den europeiska valutan under de närmaste åren .
Därför anser vi definitivt att stabilitetspakten måste iakttas bestämt och konsekvent !
Vi behöver strukturreformer inom den europeiska ekonomin .
Framför allt behöver vi en europeisk ekonomi , där det återigen lönar sig att prestera , genom att människor blir verksamma som företagare .
Det vore en olycka för Europa om det slutligen bara skulle återstå några få multinationella företag , och de små och medelstora företagen i Europa inte hade någon framtidschans !
( Applåder ) Här spelar kommissionen en viktig roll , genom att vi - tillsammans med medlemsstaterna - påbörjar en politik med skattereducering , så att företagarinitiativ återigen lönar sig .
Här vill vi gemensamt få i gång Europa .
Ni har i ert dokument talat om decentralisering och subsidiaritet .
Det stöder vi .
Nationerna , regionerna , städerna och kommunerna i Europa kommer att bevaras .
Men det finns för närvarande en utveckling - som exempel kan nämnas direktivet om livsmiljöer samt vilda djur och växter - där man åtminstone i mitt land fått det intrycket , att organisationer går vid sidan av nationella och regionala institutioner och lägger fram program i Bryssel , och att Bryssel sedan beslutar om egendom som tillhör otaliga jordbruk och företag i Europeiska unionens länder .
Jag vill bara nämna det som ett exempel på att vi måste se upp , och jag rekommenderar att man i framtiden här kommer fram till mer rättssäkerhet .
Herr kommissionsordförande , låt mig avslutningsvis säga följande : Vi har som Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater allt intresse av en stark kommission .
Om ni kan utföra ett övertygande arbete , så är det en framgång för oss alla !
Därför önskar vi er lycka till , men vi förstår vår roll också som kontrollör av kommissionen .
Om det skulle visa sig minsta tecken på att ni inte garanterar Europeiska unionens rätt - vi har för närvarande ingen anledning att kritisera detta , utan vi erkänner tvärtom att det inte ligger till på det viset - om alltså den europeiska rätten skulle kränkas , då kommer vi att bli mycket bestämda motståndare till kränkningen av denna europeiska rätt , eftersom nämligen freden i Europeiska unionen grundas på denna rätt .
Denna rätt och freden måste vi bevara i Europeiska unionen , ty det är förutsättningen för att vi också skall kunna verka som fredsstiftare i världen .
( Applåder ) Fru talman , herr kommissionsordförande !
Jag vill börja med att välkomna denna framställning av och unika debatt om regeringens - ett ord som ordförande Prodi och även jag är förtjusta i- kommissionens program för hela mandatperioden .
I första hand för att det innebär att vi kan förklara för våra medborgare vad vi har för avsikt att göra och vad vi redan håller på att göra .
Dessutom måste vi beklaga och med tanke på framtiden försöka rätta till den nuvarande situationen : det har tagit oss nästan elva månader - ordförande Prodi blev föreslagen på toppmötet i Berlin i mars i fjol - att skapa ett lagstiftningsprogram .
Felet är inte enbart hans ; vi håller på att övervinna en kris , men jag anser att det lämpligaste , med tanke på framtiden , är att tillsättandet av nästa kommission sammanfaller med framläggandet av ett lagstiftningsprogram .
Vi håller på att göra förändringar , men situationen är komplicerad .
Ordförande Prodi inledde sitt tal genom att ta upp en paradoxal situation , en paradox inom Europeiska unionen och även i världen som sådan : vi står på tröskeln till ett nytt konfessionslöst årtusende , som styrs av spindelnätet Internet och de biotekniska framgångarnas häxkonst ; faktum är att vi upplever övergången till en ny epok , men om vi begränsar oss till det som i dag är Europeiska unionen och talar om regeringar och regerande - som åtminstone på spanska för tankarna till det tidigare namnet på inrikesministeriet , men kanske är det också intressant att tala om regerande - , så är det viktigaste att Europeiska unionen får en bra regering och eftersom ordförande Prodi alltid försvarar sin födelseort Bologna , råder jag honom att åka till Siena för att ta sig en titt på något som vi alla begriper oss på , nämligen Ambrogio Lorenzettis fresker , där han skildrar bon governo och mal governo .
Det vi behöver här är en bra regering , fru talman .
Eftersom vi håller på att hämta oss efter en mycket svår kris , måste vi försöka fylla våra institutioner med innehåll och lyfta fram dessa .
Jag vill för parlamentet nämna ett faktum som vi ofta glömmer , nämligen att tillsättandet av Prodis kommission i september förra året vann starkt stöd i omröstningen , något som enligt vår uppfattning är tecken på en reformvänlig och europavänlig majoritet .
Jag vill emellertid påpeka att man i samband med denna breda överenskommelse i vissa grupper sade att majoriteten av parlamentet bör utgöra en opposition till en majoritet i rådet .
Det skulle utgöra ett hinder för något viktigt , nämligen utvecklandet av medbeslutandet i lagstiftningsprogrammet .
Jag påpekar detta , eftersom jag anser att stödet till kommissionen måste ske kontinuerligt under hela mandatperioden .
Å andra sidan får vi ta del av det politiska Europas födelse , en gemenskap med värderingar som vi delar , en europeisk union i medborgarnas tjänst .
Vad beträffar den senaste tidens händelser vill jag säga - och det kommer jag att säga den dag eller i början av den vecka som regeringskonferensen inleds - att vi verkligen måste lägga större vikt vid och lyfta fram arbetet med stadgan för de grundläggande rättigheterna som jag , efter det som vi har sagt till följd av den österrikiska krisen , absolut anser bör ingå i fördragen .
Jag tvivlar inte ett ögonblick på detta och ser det som en viktig faktor .
Därför , fru talman , vill jag även påpeka att vi måste vara medvetna om och försiktiga med vårt språkbruk .
Förra veckan beskrev den österrikiska koalitionens nya finansminister det österrikiska parlamentet som en komedi och en teater .
Vi som har tvingats leva under en diktatur vet att en diktatur kan råda med ett skuggparlament .
Däremot är det ingen demokrati utan ett levande parlament .
Jag tror att ett sådant språkbruk är extremt farligt , och fördömer härmed detta .
Vad beträffar de fyra viktigaste prioriteringar som ordförande Prodi ständigt hänvisar till , vad beträffar analysen av de utmaningar som väntar , vill jag påstå att vi är helt överens .
Jag vill ändå påpeka för kommissionen att den socialistiska gruppen har förändrat sin syn på prioriteringarna .
Vi uppfattar det som att den första prioriteringen är den ekonomiska och sociala agendan , som inbegriper det som i era prioriteringar kallas livskvalitet , det vill säga medborgarnas rättigheter som konsumenter och även som individer i förhållande till sådant som vi alltid bekräftar , men som vi inte poängterar tillräckligt , så som den europeiska sociala modellen och anpassningen av den till nya situationer , konsumenternas rättigheter samt respekten för miljön och en hållbar utveckling .
När man talar om löftet om full sysselsättning , måste utgångspunkten vara att full sysselsättning i dag inte , som på Beveridges tid i slutet av andra världskriget , enbart innebär sysselsättning för familjens manliga överhuvud .
Vi måste bekräfta jämlikheten mellan könen , den så omtalade gender mainstreaming , som är en av de punkter som är minst utvecklad i kommission Prodis program .
Det förutsätter en prioritering av jämlikheten mellan könen , en anpassning av den sociala modellen och i synnerhet en tydlig kamp mot populismen i ett läge då vår ekonomiska och sociala sammanhållning är hotad , och det bör också vara den främsta prioriteringen i kommissionens arbete .
Det bör förstärkas genom en tydlig kamp mot rasism och intolerans , så att man i praktiken bekräftar framväxten av en union som numera har en stark attraktionskraft på den övriga världen och som har förvandlats till ett område för immigration tack vare sin framgång och befolkningens höga medelålder .
Jag anser att det är det första mål vi bör uppnå .
I det sammanhanget vill jag nämna ytterligare en faktor , nämligen den ekonomiska regeringen med en gemensam valuta - jag tror att den kommer att slå igenom- och även på den punkten måste kommissionen göra framsteg .
Jag skulle vilja ha - det vill säga min grupp skulle vilja ha - en större tydlighet vad beträffar granskningen av Agenda 2000 , angående de ambitiösa målsättningarna och i synnerhet något så viktigt som kommissionen har gjort , nämligen att anamma utvidgningen i förhandlings- och integrationsprocessen .
Föreställer sig kommissionen en granskning först i slutändan ?
Frågan om beskattning betraktar vi också som en nyckelfråga .
Vad gäller regerandet i allmänhet , kan det vara intressant att göra vissa teoretiska överväganden .
En sak vill jag påpeka : det är farligt att härifrån ompröva Europeiska unionens regerande .
Jag är definitivt en anhängare av subsidiaritetsprincipen .
Om vi lyckas definiera det område vi skall regera inom , tror jag att det skulle vara mycket positivt .
För övrigt anser jag att våra överväganden även skall gälla subsidiaritetsprincipen .
Detta ska inte enbart gälla kommissionen - även våra stater , våra parlament och vårt civila samhälle måste överväga subsidiaritetsprincipen .
Slutligen , fru talman , vill jag kort hänvisa till det sista mål , som enligt vår uppfattning är högst grundläggande : en stabilisering av kontinenten och ett stärkande av Europas roll i världen .
På den punkten vill jag påstå att det råder enighet och att det finns ett stöd vad gäller prioriteringen av sydöstra Europa , utvidgningen och - det har jag redan påpekat - integrationsprocessen och stärkandet av programmet Europa-Medelhavsländerna samt av vår förmåga att förebygga konflikter , och en fråga som diskuteras mycket , nämligen utmaningen norr-söder .
Vi får inte glömma Afrika som är den kontinent som inte bara Gud utan även Europa glömde , inte heller vårt viktiga bidrag till utvecklingssamarbetet .
Och slutligen ett område på vilket vårt ansvarstagande ständigt växer , som världens främsta ekonomiska och kommersiella maktfaktor , nämligen som Europeiska unionens röst i världen , något som inte bara förutsätter en aktiv attityd inför Millennierundan .
Det förutsätter även en reform av Förenta nationerna och av de internationella finansinstituten , och där har Europa ett enormt ansvar .
Framför allt måste vi , fru talman och mina damer och herrar , kunna ge uttryck för detta i tydliga ordalag genom att i vissa avseenden ändra den jargong som vi använder oss av , för vi kan inte förvänta oss att européerna , som lever i en tid av genomgripande förändringar , skall ansluta sig till oss med entusiasm om vi fortsätter med ett internt språkbruk över deras huvuden .
Det är den främsta metoden att öka och stärka det förtroende som jag hoppas , i vilket fall som helst kommer att kunna mätas i nästa Europaval .
Kommissionens ordförande , får jag framföra till er å min grupps vägnar att vi stöder helt den utgångspunkt , kärnpunkten i analysen och den strategi som ni för fram i denna kammare i dag , nämligen att det nu obestridligen handlar om politik .
Det handlar om politik därför att vi går framåt .
Även om vi ännu inte avslutat att bygga upp alla ekonomiska system går vi vidare från den typen av funktionalistiskt byggande av Europa till ett mycket mer utmanande politiskt perspektiv .
Utvidgningen är en politisk utmaning .
Utmaningen att skapa ett område för rättsskipning och inrikesfrågor , att hantera frågor om asyl , invandring och brott är mycket politiska frågor .
Utmaningen med en gemensam utrikes- , säkerhets och försvarspolitik är en mycket politisk fråga .
På grund av att det handlar om politik är det mer komplext .
På grund av att det handlar om politik är det mer känsligt när det gäller suveränitet .
På grund av att det är mer känsligt i fråga om suveränitet är det mer känsligt när det gäller väljare och medborgare .
Vi är därför tvungna hitta en metod för hur vi skall gå vidare mot dessa politiska mål och för att ta itu med inte bara den skepsis utan den största faran , den likgiltighet som ni har identifierat .
Metoderna att åstadkomma detta är komplicerade men reella .
Jag instämmer med er åsikt att vi behöver mer synergieffekter mellan våra institutioner , inte bara mellan kommission och parlament utan också mellan dessa och rådet för att understryka den politiska utmaningens omfattning .
Vi behöver mer dialog , inte bara med varandra utan även med det civila samhället .
Vi behöver ytterligare klargöranden om vad Europatanken handlar om .
Vi måste kunna möta rädsla och oro , därför att många gånger är den största faran själva rädslan .
Med mer dialog och klargöranden kan vi kanske övervinna något av detta .
Min grupp är särskilt lockade av de kreativa möjligheter ni signalerar om utsikten om en vitbok nästa vår på området förvaltning .
När vi betraktar Europanätverket som ni beskriver är det mycket viktigt att Europa inriktas på sin kärnverksamhet , att vi har modet att föreslå områden där Europa kanske får stå åt sidan .
Det skulle kunna övertyga människor att Europa med hänsyn till förvaltningen inte är något som sköts enbart från Bryssel , som koncentrerar och drar till sig mer makt , mer beslut , mer befogenheter .
Det är den politiska kärnan i utmaningen och jag tror att ni har identifierat detta bra i denna kammare i dag .
I min grupp är utvidgningen den mest prioriterade frågan mot vilken alla andra möjligheter till reform måste mätas , antingen det gäller förvaltning , regeringskonferensen eller reformen av institutionerna .
Vi ser på utvidgningen som en partnerskapsprocess , inte som en process om " dom och oss " .
Vi ser på utvidgningen som en positiv vinst för medlems- och kandidatländer .
Jag föreslår kommissionen , som ett källa till en betydande mängd detaljerad information om utvidgningen , att lägga fram ett dokument i vilken utvidgningens betydelse klargörs , inte bara i budgetmässiga och ekonomiska termer utan i en vidare mening ; ett dokument , som Cecchinirapporten före Enhetsakten , i vilken man förklarar för människor på ett sätt som engagerar dem i debatten att detta är den stora historiska utmaning som Europa står inför i dag .
Vi måste kunna förankra dessa frågor noggrant .
Rörande den sydöstra delen av Europa håller jag med er att vi bedömer politiska institutioner efter vad de åstadkommer .
Under den tidsrymd som kommissionen och detta parlament finns till måste vi lyckas med uppgiften att uppnå den svåra och osäkra freden i sydöstra Europa .
Vi ger vårt bifall till stabiliserings- och associeringsavtal men vi skulle vilja se mer .
Vi skall offentliggöra detta material och presentera det under debatten om Swobodabetänkandet senare denna vecka .
I det strategiska dokumentet understryks Europeiska unionens globala roll .
Vårt centrala mål måste vara att ge unionen inflytande i globala frågor i proportion till dess betydelse avseende stöd , handel och finansiering .
I början av detta årtionde måste vi veta på förhand hur våra institutioner kommer att utvecklas internationellt innan nästa börjar och i synnerhet var vi passar in i internationella monetära organ , var vi passar in i FN-organ och så vidare .
Vi måste starta den debatten .
Som avslutning denna morgon , dagen efter Alla hjärtans dag , skriver tidningarna att er bröllopsresa är över .
Jag vet inte om ni är romantisk eller inte , herr Prodi .
Kanske är detta något mycket oromantiskt att säga en sådan här morgon .
Vi i den liberala gruppen välkomnar dock detta för det innebär att vi nu kan börja arbeta .
Det är som det bör vara .
Beträffande de många adjektiv ni använde i ert tal för att beskriva Europa - ett energiskt Europa , ett företagsamt Europa , ett Europa som har ett mänskligt ansikte och är vittomfattande - låt mig med ett ord som mina liberala kollegor håller mycket kärt lägga till ett adjektiv , en beskrivning av den typ av Europa vi önskar se i er strategi för förvaltningen : ett möjliggörande Europa .
( Applåder ) Fru talman , ärade kommissionsordförande !
Jag värderar högt den öppenhet med vilken ni medger att unionen i grunden måste ändras .
Ni dryftar mycket grundläggande frågor i ert program .
Jag tror att medborgarna börjar intressera sig mera för politik om vi tar fram stora frågor vid sidan av de små vardagliga ärendena .
Samtidigt måste man dock säga att ert program i många avseenden tyvärr påminner om ett partiprogram .
Det innehåller nämligen många goda avsikter men saknar i stor utsträckning konkreta förslag på hur allt detta skall genomföras .
Liksom vilket partiprogram som helst innehåller det också många inre motsättningar .
Jag skulle genom mitt eget inlägg vilja hjälpa er att identifiera dessa inre motsättningar .
För det första angående ekonomin och den sociala utvecklingen : Man måste kunna dryfta hur vi skall förena målsättningarna för konkurrens med dem för full sysselsättning ; detta omnämns ju i ert program .
Borde man när allt kommer omkring utveckla ett konvergenskriterium där man - vilket ni faktiskt antyder i detta program - ställer upp som mål att arbetslösheten inte i något medlemsland får vara högre än i låt oss säga de tre länder som lyckas bäst i den här saken ?
En ekologisk skattereform är det som min grupp vill prioritera .
Vi kan nämligen skapa sysselsättning och hållbar utveckling endast genom att ändra skattestrukturen , men tyvärr är detta - som vi alla vet - ett område där Europeiska unionen är helt oförmögen att handla .
Var vänliga och ta upp denna fråga på regeringskonferensen .
Europeiska unionen erhåller befogenheter endast genom att koncentrera sig på uppgifter som de enskilda länderna inte kan sköta på egen hand .
I det här avseendet delar säkert parlamentet er uppfattning om vikten av överstatligt beslutsfattande .
En inre motsättning i ert program berör globaliseringen .
Jag tycker det är mycket bra att ni tar upp begreppet " global kontroll " , liksom också andra här har konstaterat .
Tag dock även lärdom av händelserna i Seattle : Man måste förena å ena sidan fri världshandel och å andra sidan allt det ur mänsklig synvinkel värdefulla som vi vill värna om .
Ni måste inleda en dialog med medborgarsamhället .
Var vänliga och demokratisera de internationella organisationerna .
Europeiska unionen skulle kunna spela en avgörande roll i den process , där Förenta nationerna och Världshandelsorganisationen verkligen ställs under demokratisk kontroll .
Vi kan lägga fram motioner om detta tillsammans med er .
Slutligen ser jag det som mycket positivt att ni så ofta talar om medborgarsamhället , men detta utgör tyvärr en inre motsättning .
Ni borde också dra slutsatser vid regeringskonferensen .
Man måste ta initiativ så att medborgarna verkligen direkt kan påverka beslutsfattandet .
Det ni nyss sade oss är alldeles sant : Människorna vill ha en mera aktiv demokrati .
Detta är enligt min mening den enda möjligheten om vi vill att folk skall acceptera Europa och intressera sig för Europa .
Fru talman !
Min grupp var bland dem som ville ha ett dokument för att snarare kunna ha ett utbyte inom gruppen om kommissionens strategiska mål före debatten än att bara kunna avge en direktreaktion på ett uttalande i plenarsammanträdet .
Den främsta fördelen med texten i detta meddelande är således , enligt vår åsikt , att den finns till .
Vi är dessutom inte likgiltiga för vissa påståenden som görs i den eller avsikter som framförs , och som Prodi i sin tur just har understrukit och rent av klargjort i vissa punkter på lämpligt sätt .
Ja , den aktuella globaliseringsprocessen är , jag citerar " snarare uteslutande än inbegripande och har ökat orättvisorna " och därmed bör Europeiska unionens ambition vara att bidra till , jag citerar igen , " att nya spelregler fastställs inom unionen och i de internationella förbindelserna " .
Ja , många av våra landsmän är , jag fortsätter att citera , " modlösa och ångestfyllda " , för att de inte får se verkliga och hållbara lösningar på väsentliga eller existentiella problem såsom arbetslöshet och social uteslutning vilket påminner oss om det som bör vara en av våra absoluta prioriteringar .
Ja , vi måste tänka om i fråga om många aspekter av den aktuella gemenskapspolitiken om vi vill lyckas med det stora men svåra utvidgningsprojektet och vi behöver också , jag citerar , " ha rent strategiska partnerskap med våra grannar från söder och från öster för att bidra till stabilitet och fred " .
Vi saknar då inte områden på vilka vi kan inleda allvarliga diskussioner .
Vi kommer att noggrant granska de anmälda vitböckerna och på ett konstruktivt sätt delta i de mångtaliga påbörjade och utlovade uppbyggnadsplatserna .
Därför kommer jag nu att lämna tre kritiska synpunkter som tycks oss behöva höras om vi verkligen vill , inte bara i ord utan i sak , " utforma det nya Europa " för att använda den ambitiösa titeln på kommissionens dokument och Prodis tal .
Den första kritiska synpunkten , och i mina ögon den allvarligaste , åsyftar en viss tendens till en litet storvulen självförnöjelse från kommissionens sida när det gäller Europeiska unionen själv och en summarisk och rent av nedlåtande syn på våra partner .
En perfekt demonstration på denna frånstötande last finns i de första raderna i kommissionens meddelande .
Man talar där om Europeiska unionen såsom " ett levande bevis på att fred , stabilitet , frihet och välfärd kan ges åt en världsdel och såsom en modell för hela världen som visar den rätta vägen framåt " innan den avslutar med " att våra grannar har möjlighet att ansluta sig till denna välfärd och att vi har ett drömtillfälle för att göra det möjligt för dem " .
Jag tror att en mer nyanserad och sträng diagnostik skulle vara på sin plats .
Den idé enligt vilken euron skulle ha främjat ett samförstånd om återhållsamma löner verkar dessutom inte bekräftas av Europeiska centralbankens nervösa och upprepade ålägganden till facken , som bedöms vara alltför krävande .
Min andra kritik utgår egentligen från den första .
Denna extrema svårighet att se verkligheten i sina motsägelser och , i detta fall , att än en gång ifrågasätta sig själv ligger bakom de allvarliga begränsningar som så lägligt anges av Prodi , av viljan att bemöta medborgarnas krav .
Till exempel åtminstone vad gäller de länder som jag känner väl , tvivlar jag på att den avsikt , som upprepas tre eller fyra gånger i kommissionens dokument , att , jag citerar , " reformera systemen för social trygghet , hälsovård och pension i Europa i ett sammanhang av inbesparingar av offentliga utgifter " bemöter de personers förväntningar vars förtroende vi säger att vi vill återvinna .
Min tredje kritik är resultatet av de båda iakttagelserna : den svaga diagnosen och låsningarna på vägen till de nödvändiga förändringarna leder till ett projekt som verkar omfattas av ett svårt handikapp på grund av mångfalden av allmänna idéer , en litet impulsiv metod och därmed också av brist på uthållighet .
Men ingenting är förlorat .
Det handlar om en utgångspunkt , vi har fem år på oss för att lyckas , i den mån den politiska viljan finns och uttrycks med tillräcklig kraft och tydlighet .
Min grupp är för sin del fullt ut besluten att bidra till det .
Fru talman !
Att reformera och demokratisera Europeiska unionens institutioner är avgörande för den historiska och moraliska utmaningen om utvidgningsprocessen .
Detta var öppningsanförandet av kommissionens ordförande , Prodi , när han presenterade Europeiska kommissionens strategiska mål för de kommande fem åren .
Vi väntar på vitboken om Europeiska unionens förvaltning och avvägningen mellan medlemsstaternas regeringar och Europeiska unionens institutioner som skall offentliggöras i sommar .
I denna speciella fråga anser jag det viktigt att vi tar upp reformen av kommissionens interna beslutsprocesser .
Kommissionen har i sitt förslag till den förestående regeringskonferensen angivit att den föredrar att se mindre medlemsstater förlora sin automatiska rätt att nominera en ledamot till Europeiska kommissionen .
Detta gäller ett scenario där Europeiska unionen har över 25 medlemsstater som medlemmar .
Jag vill verkligen inte se en europeisk union byggas i två skikt .
Jag anser att detta skulle strida mot Romfördragets anda och syfte och alla andra senare fördrag .
Det måste finnas likställdhet vad gäller nationell representation inom kommissionen och inom alla andra Europeiska institutioner .
Jag vill påminna dem som strävar efter att ta bort rätten för små medlemsstater att nominera en europeisk kommissionär att USA ger små stater samma erkännande som större stater i Förenta staternas senat .
Nästan var och en av de 50 staterna i USA har två valda ledamöter i Förenta staternas senat , oavsett dess befolkningssiffra .
Varje framtida reform av Europeiska unionens fördrag kommer at kräva en folkomröstning i mitt land .
Det skulle bli mycket svårt för dem som föreslår en " ja " röst för ett sådant framtida fördrag att få stöd av det irländska folket , om vi förlorar vår rätt till vår kandidat till Europeiska kommissionen .
Otvivelaktigt skall reformeringen av Europeiska rådet också innefattas i denna vitbok om Europeiska unionens förvaltning som skall offentliggöras i sommar .
Återigen finns speciella politikområden som borde falla under de nationella medlemsstaternas ansvar .
Jag tror inte att det finns ett brett stöd i Europa för att införa kvalificerad majoritetsröstning om beskattning , rättskipning och inrikes- och utrikesfrågor på Europeiska unionens nivå .
Enligt artikel 99 i Romfördraget måste beslut fattade på EU-nivå om skatteändringar för närvarande vara enhälliga .
Jag anser att detta förslag bör kvarstå då en generell europeisk beskattningskod skulle försämra snarare än öka Europeiska unionens verksamhet .
Jag stöder utvidgningen av Europeiska unionen .
Jag stöder institutionella förändringar för att kunna garantera att utvidgningen av unionen sker på ett effektivt och strukturerat sätt .
Vi måste emellertid komma ihåg att den allmänna opinionen på 370 miljoner människor i den Europeiska unionen är en viktig faktor då man förändrar EU-fördragen .
Förändringar bör inte ske alltför snabbt och får inte vara alltför vittgående , i annat fall kommer den allmänna opinionen att göra en ratificering av varje framtida EU-fördrag mycket svår att få igenom .
Fru talman !
Jag skall tala för de radikala italienska ledamöterna .
Herr ordförande i kommissionen , ni sade nyss att inga politiska instanser upprättar femårsplaner .
Detta är sant om vi tänker på Rysslands planer på trettiotalet , men ni meddelade själv för några månader sedan , när er mandatperiod började , för talmanskonferensen att ni faktiskt skulle lägga fram ett program för mandatperioden , det vill säga de stora linjerna för den europeiska regering ni leder och vars verksamhet vi ägnar oss åt i dag .
Om det nu än skall vara ett regeringsprogram eller ett tendentiöst program ger en analys av det dokument ni har överlämnat till oss och det tal som åtföljde det inte annat än en katalog över goda avsikter eller snarare över frågor som är på tapeten , utan att man får intrycket att kommissionen tar klar ställning i någon av dessa frågor , det vill säga utför den uppgift som tillkommer Europeiska kommissionen .
I detta parlaments kammare har vi tidigare upplevt stora debatter om stora strategiska val som kommissionen har framfört , i kraft av sin initiativrätt , mer som ballon d ' essai , som förslag som sedan har rönt mer eller mindre framgång , men som ändå har bidragit till att Europeiska unionen har integrerats och utvecklats .
I detta fall har vi verkligen ett antal budord , herr ordförande : man räknar upp en hel rad frågor men ger , om ni tillåter , intrycket att kommissionen inte på någon punkt på något sätt vågar säga " i fråga om detta skulle vi behöva göra så här " .
Jag tycker bara ni verkligen tryckte - för mycket tycker jag - på en punkt , det vill säga på att den uppgift ni ser som den nästan högst prioriterade är att avveckla " onödig " verksamhet .
Låt oss emellertid se upp , herr ordförande , för vi har haft en förtroendekris för kommissionen och vi har satsat på den här kommissionen - åtminstone har en majoritet av detta parlament satsat på den här kommissionen - just för att reformeringen av kommissionen framför allt skulle innebära en förstärkning , en ny identitet , en ny medvetenhet om att åter ledas av en säker hand .
Låt oss tänka oss att kommissionen skulle vilja avveckla eller skulle erbjuda sig att avveckla till exempel de befogenheter den har fått genom fördragen , att verkställa den gemensamma politiken , eftersom den inte tyckte sig vara kapabel till detta .
Vad är det vi begär av en regering ?
Vad begär vi av denna tvetydiga och speciella så kallade struktur , Europeiska gemenskaperna ?
Det är bra att de gemensamma resurserna har en övernationell regering och att de inte delegeras till medlemsstaterna eller Kontoren för tekniskt bistånd ( BAT ) , vilket har hänt tidigare .
Ni verkar föreslå oss samma meny men på ett sämre sätt , eftersom ni som ni säger begränsar er till uppgiften att skapa någon vitbok , som ni erbjöd oss .
Det jag fruktar - även om ni skakar på huvudet , herr ordförande - är att detta betyder det som vissa länder tycker sedan många år , det vill säga att kommissionen skall vara ett bra sekretariat till ministerrådet .
Om det är denna roll kommissionen avser att spela under de kommande fem åren är vi , som är övertygade federalister , säkra på att detta inte är rätt väg att gå och vad detta beträffar kommer vi att ställa er till svars och bedöma vad kommissionen har för avsikt att göra .
Reformen är viktig men om den leder till en kantstött kommission , till att dess övernationella befogenheter reduceras och försvagas , handlar det om systemet för den europeiska integrationen , det som grundarna skapade för Europeiska kommissionen .
Vad de andra punkterna beträffar , herr ordförande , tar jag den om ekonomisk politik och socialpolitik som exempel : visst befinner sig den europeiska sociala modellen i djup kris , visst är arbetslöshetsproblemet det främsta problemet som inga av våra politiska åtgärder har lyckats lösa - och inte av en tillfällighet , men det är inte så att det kan lösas genom att man sammanställer den problemlista vi talade om tidigare , utan att ha en klar vision , ett förslag , det som gör att det finns ekonomier i vårt Europa vars takter hör till de snabbaste och som - inte av en tillfällighet - är de ekonomier som har förstått att sätta en flexibel arbetsmarknad och industri som främsta mål .
Om vi fortsätter att trassla in oss i förslag som hittills har burit mycket dålig frukt vet jag inte hur vi skulle kunna göra och vad kommissionen kan göra .
Detsamma gäller utvidgningen som självändamål , utan att den hänger samman med en mycket mer effektiv reform av Europeiska unionen och dess strukturer , med förslag som kommissionen lika gärna skulle ha kunnat framföra vid regeringskonferensen .
Herr ordförande , jag vill säga er någonting positivt , kanske tvärtemot somliga kollegers åsikt , vad beträffar det telegram ni skickade till den österrikiska regeringen .
Ert ställningstagande övertygade oss : ni gjorde rätt i att inte ytterligare isolera detta land .
Fast sedan får vi i handling se vilka de konkreta gesterna blir .
Herr ordförande , jag upprepar : det är en vision som enligt vår mening är något närsynt .
Framför allt saknas initiativ på de områden jag har tagit upp , till exempel vad gäller Balkan .
Är det möjligt att fortsätta att hålla Balkan utanför utvidgningen , utan att tycka att Kroatien , Makedonien och andra länder även de har rätt att vistas i detta gemensamma hus ?
Fru talman , herr Prodi !
Jag vill gärna berömma ert förslag om en genomgripande decentralisering av unionens verksamhet och fråga varför ni i så fall lägger fram en förteckning över lagar som är centraliserande .
Jag minns er företrädares tal för fem år sedan .
Han lovade precis som ni " mindre och bättre " , men Santer slutade med att ha levererat " mycket mer och mycket sämre " , och jag tror inte att ni heller kan leverera den utlovade varan .
Ni talar om en decentralisering , men centraliserar .
Förteckningen över lagar är ju en lång uppräkning av frågor där medborgarna förlorar inflytande och där ni , herr Prodi , tar bort detta från medborgarna t.o.m. när det gäller sociala frågor .
Ni talar om större öppenhet , men lägger fram förslag som sekretessbelägger handlingar som i dag inte är det .
Er kommission är de enda 20 personerna i EU som kan föreslå en minskad lagstiftningsmängd .
Det kan inga lokala politiker när man först har lagstiftat i Bryssel .
Lagkatalogen från kommissionen bör därför åtminstone åtföljas av en lika stor katalog över uppgifter som återsänds till medlemsstaterna och medborgarnas demokrati .
Annars växer ju lagmängden ständigt i Bryssel .
Vi har passerat 10 000 lagar och lika många lagändringar och ansökarländerna har fått 26 000 handlingar skickade till sig , som i det polska parlamentets behandling motsvarar 140 000 sidor .
Det är alldeles , alldeles , alldeles för mycket redan i dag .
Bryssel skall bestämma mindre och överlämna fler beslut till medborgarna , regionerna och medlemsstaterna , och de beslut som blir över skall endast handla om gränsöverskridande frågor som de nationella parlamenten inte längre kan besluta om på ett effektivt sätt .
Och arbetet i Bryssel skall ha en mycket högre kvalitet och ske under fullständig öppenhet , så att medborgarna åtminstone kan få litet " medkänsla " när Prodi och hans företrädare nu har tagit bort deras rätt till självbestämmande .
Till sist bara en kommentar till Dell ' Alba om vad grundarna drömde om : Läs de minnen som Jean Monnet nedtecknat .
Det han drömde om var ett litet , praktiskt sekretariat .
Det är inte det som Prodi är ordförande för i dag .
Fru talman !
I morse lade kommissionens ordförande , Prodi , fram ambitiösa mål för Europeiska unionen för de kommande fem åren , verkligen lovvärda mål , för att skapa en stark och effektiv europeisk närvaro kännbar i världen : framgång med utvidgning , klara utmaningen att sälja e-Europa och införa bättre förvaltningsprinciper .
Vi godtar att européer , i synnerhet den yngre generationen , måste ges ett brett perspektiv på var Europa kommer att befinna sig under kommande år .
Men hur skall vi lyckas när de tillgängliga resurserna är begränsade och våra institutioners trovärdighet inte är särskilt hög ?
Vi måste anpassa denna vision till verkligheten .
Här finns tre beståndsdelar som jag skulle vilja lämna som bidrag .
För det första behöver vi en framgångsrik europeisk ekonomi .
Vi måste se till att arbetslösheten fortsätter att minska i hela Europa , stärka trenden med privatisering och avreglering , uppmuntra till införande av informationsteknik och kunskap om Internet , visa att ett elektroniskt Europa är ett bra initiativ .
Men vi måste undvika att smyga tillbaka till gammalmodig reglering och kväva enskilda initiativ och företagsskapande .
Vi får inte vara rädda för globalisering , men vi måste också se till att vi förstår dess politiska effekt på nätverkssamhället .
Utan en framgångsrik europeisk ekonomi kan vi inte klara de kommande utmaningarna , framför allt inte utvidgningen .
För det andra måste vi se till att vi lagstiftar enbart när så krävs - subsidiaritet .
Göra mindre men bättre - en central politisk punkt hos den senaste kommissionen - måste vara målsättningen även för denna kommission .
Vi kommer att granska detta noggrant när vi skall utforma de årliga programmen om förslag till lagstiftning .
Bonde hade rätt när han sade att det finns denna föreställning om att göra mindre men bättre , och sedan får vi plötsligt se ett årligt program för år 2000 med 500 förslag och rekommendationer som verkar gå mot olika mål .
Vi måste bestämma vad som skall prioriteras och säkerställa att man får valuta för pengarna i vart och ett av dessa program .
Till sist måste vi se till att det blir en verklig och genuin reform av Europeiska kommissionen .
Ja , kommissionen - fördragens väktare - är avsedd att vara ett oberoende organ men det måste även vara ansvarigt inför europeiska medborgare genom vårt parlament .
Det informationsproblem som Bonde just nämnde behandlas som ett tecken på att kommissionen verkar begränsa informationen till oss , som medborgare och som parlamentariker , fastän vi har rätt till den enligt fördragen .
Kommissionen är egentligen inte i dag en europeisk regering .
Kommissionen avspeglar inte majoriteten i detta speciella parlament .
Vi i parlamentet har en stor roll att spela för att utforma förvaltningen i Europa .
Denna elektroniska förvaltning måste därför vara en lyhörd förvaltning så att vi faktiskt kan arbeta tillsammans och inse att var och en av institutionerna i Europeiska unionen har sin tillämpliga roll att spela .
Därför behöver vi trovärdighet , sammanhållning och tillförsikt om att vi genom att arbeta tillsammans kan återställa våra medborgares bild av Europeiska unionen .
Fru talman , herr kommissionsordförande !
Det har tidigare tagits många steg för att stärka Europeiska unionen , från euron till besluten om den gemensamma säkerhetspolitiken , ja även till beslutet av de 14 ledamöterna i kommissionen och av parlamentet i fråga om bildandet av den nya regeringen i Österrike .
Detta är beslut vars filosofi och principer jag helt delar .
Ändå ger jag er , herr kommissionsordförande , rätt i att det blir nödvändigt att ta många steg för att stärka EU , ty Europeiska unionen är varken tillräckligt stark för att bemästra den stora och absolut nödvändiga uppgiften med utvidgningen , eller tillräckligt stark för att tygla aktuella och potentiella rörelser som , milt sagt , har ett ambivalent och tvetydigt förhållande till de europeiska värderingarna beträffande demokrati , tolerans och integration av alla invånare på vår kontinent .
Det gäller inte bara för Österrike .
Unionen bekänner sig i Amsterdamfördraget till sina grundläggande värderingar , och EU : s institutioner bekräftade detta än en gång när den österrikiska förbundsregeringen bildades .
Dessa värderingar får emellertid bara full betydelse om de i detalj på ett begripligt sätt utgör delar av fördraget och slutligen också medger rättsanspråk för de enskilda medborgarna .
Artiklarna 6 och 7 i fördraget är nämligen inte tillräckliga om något skulle hända .
Därför måste kommissionen - det vill jag bekräfta och bestyrka - insistera på att stadgan om grundläggande rättigheter som skall utarbetas blir en del av fördraget och skapar bindande rättigheter , och att det finns en möjlighet att lämna in klagomål .
Därför måste kommissionen insistera på en kontinuerlig utbyggnad av det gemensamma området för frihet , säkerhet och rättvisa , och här är jag av motsatt åsikt jämfört med de båda föregående talarna .
Endast förnuftiga , genomförbara och humana principer för invandring och asylrätt kan sättas upp emot irrationella , förföriska och demagogiska påståenden från högern , från extremhögern .
Men , och det vill jag understryka , denna politik måste också åtföljas av en samstämmig och övertygande sysselsättningspolitik och en politik mot social utslagning , ty arbetslöshet , marginalisering och en ökande brist på jämställdhet är en optimal grogrund för antieuropeiska , nationalistiska känslor och handlande .
I detta sammanhang , herr kommissionsordförande , vill jag också gå in på de problem med globaliseringen som ni nämnde , och på hur stora delar av befolkningen ser på den .
Känslan av att vara utlämnad , bristande möjligheter till inflytande och bristande skydd från statens sida leder i bästa fall till att man vänder sig bort från politiken och avstår från att rösta i valet , så som skedde vid Europavalen , och i sämsta fall väljer ett extremistiskt valbeteende .
Här har unionen , vi alla , ännu inte förstått att erbjuda våra EU-medborgare EU som ett medel , ja som ett skydd mot de negativa effekterna av globaliseringen .
Vi håller på att bygga ett hus , men alltför få av våra egna medborgare känner sig verkligen hemma i detta hus .
Därför handlar det inte bara om en reform av Världshandelsorganisationen och den ekonomiska arkitekturen - och kommissionsordföranden har betecknande nog glömt bort att tala om reformen av den internationella ekonomiska arkitekturen - utan det handlar också om förtroendeskapande åtgärder för våra medborgare , som har all rätt att förvänta sig hjälp och stöd av och i EU i de oundvikliga , men smärtsamma processerna med att anpassa sig till de nya globala förhållandena .
I detta sammanhang är det som kommissionen säger om Europas styrkande röst betydelsefullt .
Ni själv , herr ordförande , har i dag talat om en modell , som jag tyvärr finner alltför litet om i dokumentet ; ni sade att vi både i inrikes och utrikes frågor måste erbjuda våra medborgare en modell för ekonomisk , social , kulturell och ekologisk utveckling , som tydligt skiljer sig från andra modeller , även från USA : s modell .
Här är USA inte heller enbart vår partner , utan också vår konkurrent , och vi måste kämpa om vem som erbjuder den bästa modellen för våra medborgare .
Jag skulle önska mig att det som vi i dag har sagt med sådan intensitet också i högre utsträckning skulle återfinnas i kommissionens dokument .
( Applåder ) Fru talman !
Kommissionens ordförande !
Den största gåvan som er kommission kan lämna över till Europeiska unionen skulle vara att medverka till en omflyttning och omfördelning av kommissionens alltmer röriga och hoprörda befogenheter och behörigheter och eventuellt för själva unionen .
Ni har gjort en djärv start genom att rätteligen understryka nödvändigheten att fokusera på de så kallade " huvuduppgifterna " .
Det innebär som ni själv framförde i dag att man också måste identifiera de arbetsuppgifter , politikområden och program som ligger utanför eller inte hör till kommissionens centrala ansvarsområden .
Många av Europeiska unionens nuvarande politikområden och program kanske helt enkelt har passerat sitt sista användningsdatum eller har befunnits vara ohanterliga eller ineffektiva när de administreras på europeisk nivå .
Utmaningen nu är att ha modet att flytta tillbaka så mycket icke-kärnverksamhet som möjligt till lägre nivåer på nationell , regional och lokal ledningsnivå .
Om vi skall lyckas övertyga en skeptisk europeisk allmänhet om fördelarna med ytterligare europeisk integrering , måste vi kunna visa att vi är lika duktiga på att fördela omotiverade befogenheter som vi är på att skapa nya befogenheter för EU .
Vi får inte låta kritikerna av europeisk integration hävda , som de för närvarande gör med visst berättigande enligt vad vi just har hört av Bonde , att ökningen av EU : s ansvarsområden endast går åt ett håll .
Det måste ses som en tvåvägsprocess där befintlig EU-politik och EU-program som inte klart kan försvaras enligt principerna subsidiaritet och proportionalitet överflyttas och avskaffas .
Om ni kan hitta åtgärder som är i linje med dessa strävanden under de kommande åren kommer ni att lämna ett exempellöst bidrag till hela Europeiska unionens framtid , och som vi har hört i dag kommer ni att få ett betydande stöd i detta Europaparlament .
( Applåder ) Fru talman , herr kommissionsordförande !
Jag samtycker fullt ut med tankarna i de förslag som gjorts av min kollega Heidi Hautala vad gäller kommissionens strategiska mål för de kommande fem åren .
Jag kommer för min del att hålla mig till ett ämne som ni inte har tagit upp och som hade planerats och gäller kommissionens arbetsprogram för år 2000 .
Jag är medveten om budgetårets begränsningar eftersom vi arbetar inom ramen för det aktuella fördraget och är begränsade av dess funktionsregler - jag tänker särskilt på en viktig fråga som är skattefrågor .
Men jag skulle faktiskt inte vilja tala om skattefrågor .
Jag kommer att börja med att välkomna vissa förslag som ni lägger fram inför programmet för år 2000 .
Jag tänker på alla förslag i fråga om livsmedelssäkerhet som är ambitiösa och viktiga och jag tänker också på sjösäkerhet efter de båda oljeutsläppen utanför Bretagnes kust och i Turkiet .
Det är bra att kommissionen reagerar snabbt i det avseendet .
När det gäller andra frågor anser jag däremot att man skulle kunna vara mer ambitiös och gå snabbare .
Och jag skulle vilja lämna ett antal positiva förslag , där tänker jag framför allt på det sociala området , miljön och uppföljningen av Seattle .
En inledande anmärkning : ni sade att det är nödvändigt att åter försona de europeiska medborgarna med deras institutioner , något som är självklart , och jag tror således att det är viktigt att vi undrar över vad som i främsta ledet upptar medborgarnas tankar .
Jag tror till exempel att på det sociala området räcker det inte med att utfärda ett meddelande om ett program för sociala åtgärder .
Det måste gå snabbare .
Ni måste lägga fram ett nytt program för sociala åtgärder för oss i slutet av året .
En fråga , slutligen , som har ingått i de senaste nyheterna och fortfarande upptar en stor plats i dem är frågan om företagsnedläggning och kollektiva uppsägningar .
Vi arbetar på grundval av ett aktuellt direktiv som har visat sig ha sina begränsningar och vi skulle vilja - och jag ger er ett förslag - se över denna direktivtext så att vi får ett effektivare direktiv vad gäller sysselsättningsskydd och också effektivare vad gäller eventuella sanktioner mot dem som inte följer texten .
När det gäller miljön aviserar ni ett förslag till beslut om ett sjätte åtgärdsprogram om miljö och det är mycket bra .
Man har sagt mig - men ni skall kanske dementera mina uttalanden - att det inte finns några exakta mål och någon tidsplan för genomförande i den text som ni skall föreslå oss .
Jag tror personligen att det är nödvändigt att ha beräknade mål och en verklig tidsplan för genomförande .
Jag tror också att när det gäller frågan om enskilt ansvar är det glädjande att vi äntligen har en vitbok , jag talar då om enskilt ansvar gentemot miljön , men jag vill påminna om att parlamentet har begärt ett lagstiftningsinitiativ i sex år , och att vitboken naturligtvis aviserar en sådan lagstiftning , men när ?
Där vill jag också uppmärksamma er på att processen måste påskyndas .
Slutligen den sista delen , efter Kyoto skulle det ändå vara sunt om vi skulle snabbt komma fram till exakta förslag och jag vill sluta med att säga ett ord om WTO .
Jag tror att tanken på att åter sätta i gång en ny global period inte är en dålig tanke men jag tror och upprepar att först måste verkligen kommissionen ge oss förslag för att ändra WTO : s funktionsregler .
Kommissionen har en inre roll , men också en roll i världen .
Det verkar som om Europeiska unionen bör ligga till grund för en omvärdering av WTO : s funktionssätt , en omvärdering som bör leda till att vi ger exakta förslag i stadgehänseende .
Fru talman !
Ni talade om grundläggande politiska värderingar och en av de grundläggande politiska värderingarna , till och med mer grundläggande än demokratin , är respekten för andra .
Därför anser vi att ni gjorde rätt i att skicka ett meddelande , och att de som kritiserar det kanske fortfarande lider av sviterna av en bolsjevitisk eller nazistisk kultur , för demokrati innebär att föra en dialog med andra och låta dem förstå när de felar , men också lyssna på deras skäl .
Att utvidga får inte innebära att urvattna , det vill säga det får inte innebära att man utvidgar riskerna .
Detta har Nationella alliansen upprepat i tio år i denna kammare .
Kandidatländernas förhoppningar är minst lika viktiga som våra nuvarande medborgares förhoppningar , vilka börjar bli allvarligt besvikna på hur detta Europa fungerar när man inte löser de viktigaste problemen .
Utvidgningen kräver alltså stränghet , att man respekterar de villkor som - om det blir nödvändigt - bör omformuleras vad vissa grundläggande frågor beträffar : det som har hänt i Rumänien , med konsekvenser ända till Belgrad - den ekologiska tragedin - men framför allt att likgiltigheten inför de stora säkerhetsproblemen fortsätter att breda ut sig .
Än i dag finns inga slutgiltiga lösningar för kontroll över kärnkraftverken i östrepublikerna .
Man måste alltså ha resurser att spendera innan man går vidare mot en utvidgning , för att äntligen skapa en europeisk kontrollstyrka med uppgift att övervaka kvalitet och driftsförhållanden för att skapa en ny värld där vissa tragedier inte längre hör hemma .
Jag skulle också vilja säga några ord om Afrika , fru talman .
Den tredje och fjärde världen är övergivna : det skulle räcka med en dollar , en och en halv euro , för att rädda många barn .
Europa som är så demokratiskt , som är så progressivt , tiger och tar inte på sig dessa tragiska problem , under tiden som halva Afrika dör i aids och andra sjukdomar .
Ett sista påpekande om Internet och globaliseringen .
Globaliseringen av ekonomin får inte bli en likriktning av produkter och kvaliteter , liksom globaliseringen av politiken inte får bli en utslätning av värderingar , av förhoppningar , av entusiasmen .
De folk som inte deltar , och som sakta drar sig undan , ger utrymme för en oligarki som tar makten och lämnar kontrollen till ett fåtal .
Vad Internet beträffar : Europa måste äntligen ha modet att säga att det krävs regler .
Tillåt mig här att , som privatperson , applådera de pirater som genom att handla som de gör tvingar världen att fundera över det enda system som inte har några regler i dag .
Vi är en reglernas värld : låt oss ge även Internet regler och på så sätt ge medborgarnas framtid regler och hopp .
Fru talman !
Som skattebetalare i Padanien har jag redan känt av uttaxeraren Prodis bett på den tiden då han var regeringschef i Italien som Padanien också skattemässigt är underställt .
Jag blev bekymrad när jag lyssnade på honom nu när han antydde nya resurser , ett koncept som lätt kan översättas med nya skatter och pålagor bland annat inför utvidgningen , det vill säga att nya stater träder in i unionen .
Men varför betalar inte de sin inträdesbiljett själva ?
Mina padanska väljare som tack vare Prodi redan har betalat det som i Italien går under namnet Europaskatt - som bara delvis har återbetalats - har absolut inte för avsikt att , fortfarande tack vare Prodi , betala en skatt till för någon annan .
Fru talman , herr kommissionsordförande , ledamöter av kommissionen !
Fem månader efter sitt tillträde har kommissionen angivit i vilken riktning den vill styra Europeiska unionen .
Det har blivit en ambitiös men även högtravande handling .
Är det inte patetiskt att säga att " världen ser upp till Europa " ?
Dessutom är världsdelen Europa så mycket mer än de femton medlemsstaterna i Europeiska unionen .
Garanterandet av fred , demokrati och mänskliga rättigheter i , märk väl , hela Europa är att sikta litet väl högt .
Jag är väldigt nyfiken på hur kommissionen tänker förverkliga det här .
Den europeiska integrationsmodellen som en rik källa för världsstyre , är det detsamma som export av storskalighet och maktkoncentration ?
Kommissionen anser att utrikespolitiken kan lyckas om var och en vet exakt vem som styr !
Vem är det då ?
Hela kommissionen , dess ordförande kanske , rådet ?
För den nya ledningen av Europa behövs starka institutioner , säger ni , medan kommissionen samtidigt vill koncentrera sig på sina kärnuppgifter .
Det senare håller vi gärna med om .
Det är verkligen hög tid att institutionerna inskränker sig till problem som verkligen är gränsöverskridande och slutar smycka den europeiska vagnen med befogenheter som tagits från de nationella myndigheterna .
Vid flera tillfällen i texten talas det om gemensamma värden .
Tyvärr saknar jag en hänvisning till de normer som hör dit .
Man kan undra var de normerna och värdena är hämtade från .
Jag är övertygad om att Bibeln , Guds ord , är den enda rena källan till goda normer och äkta värden .
Den insikten är en viktig del av traditionen i vår världsdel och den förtjänar att bli erkänd Fru talman !
Jag skulle vilja gratulera Prodi och kommissionen till deras regeringsförklaring .
Huvuddragen i den tilltalar mig verkligen .
Jag delar också Prodis och kommissionens analys att det inom flera områden finns ett behov av mer Europa , mer integrering .
För områden som säkerhet , Världshandelskonferensen , livsmedelssäkerhet och även den nya ekonomin krävs det alltså fler åtgärder av Europeiska kommissionen .
Utmaningen kommer att vara hur medlemsstaterna , rådet , Europaparlamentet , de nationella parlamenten , kommissionen och diverse andra aktörer skall kunna föras samman på en och samma linje .
Europeiska kommissionen måste i det avseendet spela en viktig roll som regissör men för det krävs tydliga och genomförbara målsättningar .
Klara prioriteter , fokus och främst även kommunikation med samhället om vad vi håller på med .
Det är de nyckelåtgärder det handlar om och för det krävs av kommissionen , med tanke på subsidiariteten , konkreta arbetsresultat som vi sedan gärna vill se i de kommande programmen .
Att tyngdpunkten läggs på kärnfunktionerna är i sig alldeles utmärkt och att kommissionen ser sig själv i en bättre , större roll med avseende på politiska koncept och politiska initiativ , det välkomnar jag .
Men vad det också handlar om , är genomförande , att verkställa det som kommissionen planerar .
Om jag till exempel ser på telekommunikationssektorn så ser jag att vi utfärdat väldigt många direktiv , men att det ändå fortfarande finns femton delmarknader och att femton medlemsstater fortfarande genomför direktiven på olika sätt .
När det då gäller genomförandet : det handlar naturligtvis också om att kommissionen ser till att det som vi vill i politiken även märks i praktiken .
När det gäller utrikespolitiken , fru talman , så är jag väldigt tilltalad av ambitionen att Europeiska unionen måste ha lika mycket politisk och ekonomisk vikt .
Jag undrar bara : när det talas om en verkligt gemensam politik , om ett system för krisförebyggande och krishantering på gemenskapsnivå , var finns de konkreta förslagen ?
Det är ju så vi måste pröva om vi verkligen kan förverkliga vår målsättning på det området .
Prodi ägnade med all rätt mycket uppmärksamhet åt Afrika i sitt anförande men jag måste säga att jag ändå är besviken när jag tittar på arbetsprogrammet för år 2000 .
Där hittar jag överhuvudtaget inga åtgärder som berör Afrika , varken i inledningen eller i själva programmet , och jag hoppas alltså att Prodi skall lägga fram ett bra meddelande som förberedelse inför toppmötet i Afrika .
Fru talman !
Ord är mycket viktiga men vi kan endast bedöma kommissionen efter dess gärningar .
Fru talman , herr kommissionsordförande , mina damer och herrar !
Jag vet inte vad jag skall hålla mig till - de strategiska målen för perioden 2000-2005 eller till ert tal om perioden 2000-2010 ?
Har ni redan inkluderat er andra mandatperiod ?
Men , allvarligt talat .
Unionen som håller på att utvidgas behöver stärkas genom bantning och begränsning .
För det första , bantningen .
Det ni säger i ert program om att koncentrera sig på kommissionens kärnfrågor är bara en första början .
Hela unionens verksamhet måste föras tillbaka till politikens kärnområden .
De omfattar marknadens sociala och ekologiska inriktning , säkrandet av valutan , garantin för de medborgerliga rättigheterna inom unionen och företrädandet av de gemensamma intressena utåt .
Här gäller det inte bara att tala med en röst i världen , utan det handlar snarare om vad vi vill säga med denna röst .
För det andra heter det nya modeordet flexibilitet .
Men en tilltagande flexibilisering kan bli eller hotar mycket snabbt att bli till ett samarbete på regeringsnivå .
Vi måste benhårt hålla fast vid sammanhållningen av medlemsstaterna med hjälp av gemensamma beslutsorgan .
Det gäller för övrigt också för införlivandet av det civila samhället , som kan betraktas som positiv .
Men medborgarna behöver inga nya organ eller institutioner och absolut inte någon ny sammanblandning av ansvarsområden .
( Applåder ) Öppenhet betyder inte större tillgång till mer papper , utan öppenhet för medborgarna är att äntligen få mer klarhet om vem som beslutar när och med vilket berättigande i Bryssel och Strasbourg .
Det är öppenhet !
För det tredje kan och får Europeiska unionen inte utvidgas gränslöst .
Dess gränser bestäms inte av hur många stater som vill vara med , utan av hur många stater som den klarar av .
( Applåder ) Om priset för utvidgningen vore en uppmjukning eller rent av en upplösning av den befintliga unionen , då får man inte betala det priset .
Det skulle vara för högt , för övrigt inte bara för dess medlemsstater , utan också för de stater som vill bli medlemmar i unionen .
En union enbart som ett geostrategiskt koncept har inte någon framtid , lika litet som en union som enbart är en frihandelszon .
Men unionen förblir något mer än en marknad och får sin legitimitet av Europas folk enbart om den uppfattar sig som en ödesgemenskap .
Detta är långt mer än enbart er nya ekonomiska och socialpolitiska agenda eller en ny och bättre livskvalitet .
Inte bara kommissionen , inte bara Europaparlamentet , utan också folken och staterna i vår Europeiska union måste finna nya svar på frågan hur och för vad vi vill leva och agera gemensamt .
Här handlar det inte om något mindre än att uppfinna Europeiska unionen på nytt , utan att förstöra det som redan existerar !
( Applåder ) Herr talman !
Enligt Europeiska liberala och demokratiska partiets grupp är kommissionens och hela unionens viktigaste uppgift under de närmaste åren att genomföra utvidgningen med framgång .
Kommissionen skall i förhandlingarna målmedvetet sträva efter att varje ansökarland skall kunna gå med i unionen snarast möjligt .
Å andra sidan måste man se till att inte omintetgöra hittills uppnådda resultat eller målsättningarna för integrationen .
För att undvika detta har den liberala gruppen framfört ett önskemål om att man vid regeringskonferensen skall överväga olika modeller för en differentierad integrering och att man skapar en koncentrisk union med en federationskärna och en mindre integrerad yttre cirkel .
Det är uppenbart att unionens interna differentiering tas upp på regeringskonferensen .
Behandlingen av denna fråga kräver fördomsfrihet .
Det räcker inte med att tekniskt förbättra det flexibla samarbetet , utan man måste också diskutera utvecklingen av de egna institutionerna för avant garde-länderna , såsom bland annat Jacques Delors har föreslagit .
På detta sätt kan vi skapa en ännu effektivare , tydligare och mera demokratisk beslutsprocess .
Jag hoppas att komissionen lämnar ett eget förslag till hur den institutionella och övriga differentieringen i den utvidgande unionen bör genomföras .
Fru talman , herr kommissionsordförande , mina damer och herrar !
Ert inspirerande anförande , herr Prodi , har förfört mig .
Det väcker förväntningar men det kan också leda till besvikelse .
Det har att göra med det som Van Velzen sade alldeles nyss , med skillnaden mellan ord och handling .
Unionens utvidgning kommer sig av vår längtan efter fred , säkerhet och stabilitet .
Ni vill lugna de nya staterna och även den europeiska opinionen .
Vi ser dock med våra egna ögon att det motsatta sker i dag .
Vi ser hur rädslan och oron ökar , även i de områden där arbetslösheten inte är hög och välfärden är väldigt stor .
Vi måste kunna ge våra medborgare en hemkänsla , sade Swoboda , och det har han rätt i .
Det är en plats där vi alla delar samma värden och där var och en har sin uppgift och sitt ansvar .
Det har antagligen att göra med de normer som Van Dam talade om .
Det är nämligen subsidiaritet .
Tydligt ansvar för alla ledningsnivåer , partner och inte konkurrenter i styret .
Makten så nära medborgarna som möjligt , där den kan utövas öppet och under insyn och kontrolleras av medborgarna själva .
För det krävs en ny politisk kultur , inte bara i teorin utan även i praktiken , där man tar hänsyn till den verklighet som råder i medlemsstaterna och i regionerna .
Regioner som i kulturellt och ekonomiskt avseende ibland är lika viktiga som vissa medlemsstaters intressen .
Det nya Europa får inte bara utvecklas på bredden utan även på djupet , genom att omsätta våra värden i praktiken och genom ett demokratiskt byggande av en äkta gemenskap .
På det skall kommissionen bedömas .
Fru talman , kommissionen lägger idag fram sina strategiska målsättningar för perioden 2000-2005 i form av ett extremt allmänt hållet dokument i vilket de sträva anmärkningarna strukits för att inte alltför mycket såra en del personer .
I den första delen således rörande de nya formerna av europeiskt regerande läser man inte någonstans naturligtvis orden federalism eller superstat .
Men det är ändå de som framträder när det är fråga om en stark europeisk institution i vilken enbart de löpande genomförandeverksamheterna decentraliseras och skjuter in sin kollektiva syn i en oklar enhet där regeringar och nationella parlament är beblandade med regionala , och till och med lokala , myndigheter samt med det civila samhället , samtliga utsedda , utan någon hierarkisering såsom , jag citerar : " deltagande part i europeiska frågor " .
Dessa tvetydigheter döljer många missuppfattningar och främst om våra värderingar .
Det räcker nämligen inte med att åberopa demokrati för att vara demokrat .
Man måste framför allt acceptera att medborgarna fritt fattar beslut på den nivå där de objektiva villkoren för en nära , lojal och öppen demokratisk debatt bäst finns samlade , det vill säga huvudsakligen på nationell nivå .
Kommissionens meddelande i sin helhet är emellertid just uppbyggt på motsatt påstående enligt vilket det skulle vara nödvändigt att under förevändning att bättre försvara folket fortsätta att begränsa deras marginal för självständigt val ytterligare genom nya föreskrifter , nytt införlivande av politik eller nya tvingande rättsliga strukturer såsom förslaget till stadga om så , felaktigt , kallade grundläggande rättigheter .
Jag betonar " felaktigt " eftersom den i själva verket skall minska dessa rättigheter .
I Gruppen Unionen för nationernas Europa är principerna mycket annorlunda .
Vi vill försvara Europas länder men också respektera folkens val .
Det är inte alls cirkelns fyrkant .
Vi måste nämligen överge de omoderna federalistiska modellerna , de modeller som satts upp av dem vars idéer om Europafrågan härrör från Jean Monnets memoarer .
Vi måste tvärtom öppna de europeiska institutionerna för den moderna världen genom att uppfinna en dynamik av variabel geometri som respekterar nationerna .
Detta är den stora idén om ett nytt ledningssätt som vi skulle ha velat finna i ert meddelande , herr ordförande .
Tyvärr fanns det inte där .
Fru talman , herr kommissionsordförande !
Ni påstår att ni utformar ett nytt Europa men ni saknar tyvärr en väsentlig förutsättning : förtroende .
Man kan nämligen inte dra till sig miljoner européers förtroende när man inte är värd det .
Och hur skulle ni kunna vara värd ett förtroende efter galna ko-affären och Santer-kommissionens avgång på grund av korruption ?
Ni bär ansvaret för miljoner arbetslösa och miljoner fattiga samt ökande utsatthet och nöd på grund av er extrema handelsutbytespolitik och ultraliberala politik och på grund av tvångsmarschen till den gemensamma valutan .
Ni har velat ha och har ordnat avlägsnandet av de inre gränserna och ni har sålunda utsatt Europa för en explosion av kriminalitet och osäkerhet och en flodvåg av okontrollerad invandring .
Ni föreslår nu att en handfull tjänstemän skall få hela beslutandemakten och göra staterna , de lokala myndigheterna och de icke-statliga organisationerna , där alla för övrigt har lika villkor i sitt beroende till Bryssel , till enkla verkställare av beslut som kommer ovanifrån .
I ert fjortonsidiga dokument nämns inte en enda gång de nationella parlamenten , som likväl i motsats till kommissionen består av folkvalda ledamöter .
Men de har visserligen inte någon roll i er strategi .
Ni vågar inte ens kalla saker och ting med sitt rätta namn och ni gömmer er bakom en låtsad inne-semantik genom att kalla det för " guvenörskap " , det som inte är något annat än en federal enväldig centralregering .
Efter att i åratal ha försökt övertyga genom att tala om delad suveränitet medger ni nu ert yttersta mål : att sälja ut den europeiska suveräniteten , vare sig den är nationell eller lokal , till en världsregering i vilken ni inte ens hoppas på att få en avgörande plats .
Ni vågar slutligen fördöma och sanktionera , eller låta fördöma och sanktionera , miljoner österrikares fria och demokratiska val av det skälet att ni inte tycker om resultatet .
Och på samma gång stöder ni det kommunistiska Kina och har handel med länder som öppet bryter mot mänskliga rättigheter sedan årtionden tillbaka .
I dag igen går de europeiska parlamentsledamöterna angrepp mot ett telegram från Prodi till kansler Schüssel som likväl påtagligen inte är en sympatiyttring utan en politisk manöver .
Ert skryt bedrar inte någon eftersom , och det vet ni mycket väl , vare sig ni vill eller inte behöver ni Österrike för att reformera fördragen och harmonisera skattesystemet för sparande .
Ni använder Österrike som en bekväm fågelskrämma .
Era kommissionärer är förvisso inte de enda som är ansvariga .
De regeringar som stöder er av slapphet eller av ideologiska skäl är det också .
Bryssel är inte vi alla som ni påstår , utan det är ni alla .
Ljug inte mer , ni struntar väl i vad Europas folk vill .
Européerna är bara fria att välja mellan er bästa av världar och att ställas vid skampålen .
Mer än tio år efter Sovjetunionens upplösning osar era förslag av gulag med tillägg av en lenande moralism .
Vi var en del av den lilla klick som pekade ut den kommunistiska diktaturen .
Vi är och kommer att förbli bland dem som bekämpar en europeistisk diktatur och vi uppmanar alla Europas folk att gå med i motståndet mot era ohyggliga förslag .
De europeiska demokratiernas räddning finns i staten såsom nation och i den nationella staten och Europas räddning finns i samarbetet mellan nationerna i Europa .
( Några applåder ) Ordförande Prodi , ni har i dag presenterat ett femårsprogram för kommissionen med många mål som man kan instämma i , ett program som består av scenarier och ledmotiv , och det är därför riktigt att hålla sig kvar vid de stora dragen , bortom de konkreta inslagen .
Av era ord och det dokument ni har överlämnat till oss verkar det som om en fråga som ligger er , herr ordförande , och mig varmt om hjärtat har hamnat i skymundan : solidariteten , inte så mycket på det internationella planet som internt .
Ärkebiskopen i Milano , Hans Högvärdighet Carlo Maria Martini , uppmanar alla politiker och särskilt sådana som ni och jag , herr ordförande , sådana som kulturellt och värdemässigt grundar sitt politiska engagemang på katolicismen , att omvärdera en utvecklingsfråga som förutom den ekonomiska vinsten mycket , oerhört mycket , berör dem som har det sämst ställt , de utstötta .
Det är en stor fråga , den om de som har det sämst ställt , en stor fråga som påminner oss om hur svårt och komplicerat det är att fastställa mått på framsteg och hur otillräckligt det är att bara se till inkomsten per capita .
Det påminner oss också om behovet av en ny utvecklingsmodell som är stadigt förankrad i en kultur med socialt engagerade katoliker , vilka betraktar det civila samhället , de samhälleliga instanser som allmänheten främjar och understöder , som de sundaste instrumenten för att bygga solidaritet .
På så sätt betonas den grundläggande elementet för varje individs utveckling : hennes frihet , som kommer före den ekonomiska vinsten .
Denna samhälleliga frihet som yttrar sig i initiativ till förmån för dem som har det sämst ställt ger återbetalning i form av rättvisa och samhällelig balans .
Herr ordförande , de offentliga institutionerna skall inte bara följa ekonomiska kriterier .
De måste rikta in sig på service till individerna och arbetet med att bygga upp var och ens frihet , naturligtvis utan att glömma att allt detta inte får och inte skall stå i motsats till behovet av att skapa företagsamhet , att investera och riskera .
I ett ordentligt och målinriktat system kan entreprenörerna bidra till samhällets tillväxt och till solidariteten i betydande omfattning .
I globaliseringens tidevarv , globaliseringen som vi dock vill ge en ram av fasta regler som ger de ekonomiska aktörerna och konsumenterna trygghet , får inte Europeiska kommissionen glömma solidariteten och betona att den skall tillämpas i alla medmänskliga relationer .
Vår historia har lärt oss att hjärtat måste finnas med i politiken .
Vi hoppas att vitboken och era och kommissionens handlingar kommer att visa detta i praktiken .
Fru talman , kommissionsordförande , kolleger !
Shaping the new Europe är en ambitiös målsättning för kommissionen och för oss alla .
Vår ambition och vårt arbete kommer att följas av medborgarna i våra länder , men också av många utanför Europa och utanför vår union .
Vilken bild får då en intresserad allmänhet och resten av världen av detta femårsprogram ?
Mitt svar är : en nystart , en tydligt reformistisk agenda , som bekräftar att 2000-talets union inte vill stanna vid att vara en ekonomisk gemenskap , utan vill vara en värdig gemenskap , som vi tar på allvar .
Med rätta säger kommissionen att unionens avsikt är att utveckla och värna om ett solidariskt välfärdssamhälle i globaliseringens tidevarv , ett rättfärdigt och effektivare Europa , som också ser sitt ansvar utanför den egna kontinenten utifrån solidaritet och upplyst egenintresse .
Vi ser nämligen fattigdom och utanförskap som fredens och frihetens främsta fiende .
Med instämmande i vad mina partivänner har sagt och med gillande av grundtonen i ert dokument vill jag rikta uppmärksamheten på två brister , som måste korrigeras i det kommande arbetet .
Det första gäller kvinnor , gender eller kvinnors rättigheter .
Ni talade om kvinnors medverkan för att öka produktion och tillväxt .
Detta är viktigt , men jämställdhet är inte bara nödvändigt för produktiviteten utan också för demokratin i våra samhällen .
Det är därför uppseendeväckande att ordet jämställdhet , gender eller kvinna överhuvudtaget inte förekommer någonstans i Shaping the new Europe .
Ni talade om kvinnan i ert tal , men hon nämns inte bland de strategiska målen .
Beror detta , herr kommissionär , på att mainstreaming redan är så genomförd i kommissionen att kvinnor inte behöver nämnas ?
Hur förklarar ni annars denna frånvaro av kvinnor .
EU får inte bli en union med manligt ansikte .
Min andra fråga gäller Afrika .
Inte heller Afrika nämns i Shaping the new Europe , men alla andra kontinenter .
I Afrika har vi världens högsta antal flyktingar , världens största samlade fattigdom och en förtärande aidsepidemi .
Jag vet att kommissionär Nielson och andra gör ett bra jobb , men det krävs att hela kommissionen , också i sina strategiska målsättningar , fokuserar mer på denna kontinent .
Slutligen vill jag välkomna kommissionens uttalande och att det i detta för första gången sägs att EU är berett att unilateralt vidta åtgärder till förmån för ökat tillträde till våra marknader för utvecklingsländerna .
Min fråga är : När kommer detta att sjösättas ?
Fru talman , herr ordförande i kommissionen , ärade ledamöter !
Vi har framför oss ett dokument som har avgörande betydelse för Europas framtid och öde .
Av alla frågorna framträder emellertid direkt två som är intimt förknippade med varandra : freden och stabiliteten i och utanför Europa .
Det handlar om mål som skall prioriteras .
Sedan länge delar vi alla detta synsätt , men vi måste också tydligt hävda att dessa mål inte kan uppnås utan utvidgningen , även om denna skulle medföra kostnader .
I dag är det vår uppgift att för de kommande decennierna välja mellan ett Europa som kanske är mindre rikt , men som är en ledstjärna för fred och civilisation för hela vår planet och ett Europa som kanske är mer välmående men saknar visioner .
Dessa mål kan dock endast uppnås om regeringskonferensen , som kommer att avslutas innan årets slut , ger upphov till en konstitutionell reform som ger kommissionen adekvat och reell makt .
Kommissionen kan inte fortsätta att bara vara den som verkställer rådets beslut och parlamentets medbeslutande utan måste spela rollen som Europas verkliga regering .
Parlamentet borde vara den förste att stödja denna reform om det verkligen vill vidga sin roll som uttolkare av européernas vilja och skaffa sig den centrala funktion som tillkommer en union som är sant demokratisk och kraftigt integrerad .
För övrigt kan kommissionen bara ges ansvar för de åtaganden den tar på sig i den utsträckning den reella befogenhet den har medger .
Om dessa skisserade möjligheter saknas kommer Europa att retirera in i en historia utan framtid .
Fru talman , herr kommissionsordförande !
Vi kan glädjas åt den globala ambitionen i de angivna målsättningarna , som går parallellt med de utmaningar som Europa skall tvingas klara av .
Jag noterar att ni anser att Berlinmurens fall är den väsentliga faktorn i sekelslutet .
Denna händelse bör leda till utvidgning .
Jag har lust att snarare tala om återförening än att använda ordet " utvidgning " .
Det tycks mig ha en politiskt mycket starkare betydelse .
Ni återupptar tanken att omcentrera era verksamheter runt de viktigaste uppgifterna och det ingår i målsättningarna för er reform .
I grunden handlar det om att tillämpa subsidiaritetsprincipen .
En klar tillämpning av denna princip kan bara stärka de åtgärder som vidtas och ge medborgarna en klar bild av varje behörighetsnivå .
Men , herr Prodi , att säga det är en sak men att göra det är en annan !
Ni måste således kämpa mot alla institutioners tendens att i allmänhet försöka öka sina befogenheter ytterligare .
Jag kommer således att döma efter handling .
Under tiden instämmer jag i och uppmuntrar denna tydligt uttryckta vilja i ert meddelande .
Två saker är emellertid väsentliga : förenkling och tillämpning av gemenskapsrätten .
1998 var det 123 anhängiggöranden i domstolen på grund av icke-tillämpning eller icke-införlivande av gemenskapsrätten och 25 procent av direktiven om miljöfrågor tillämpas inte eller är inte införlivade .
Händelserna de senaste dagarna visar hur nödvändigt det är .
Gemenskapsrätten får inte vara utan tillämpning för att den är för komplicerad eller för detaljerad .
Unionen får inte falla i den fällan och också i det avseendet beklagar jag att ert meddelande inte går in mer på detaljer .
Ni är realistisk i fråga om att välfärdsstaten inte längre kan lösa de problem som uppstår och bland annat arbetslösheten .
Jag beklagar dock att ett klart alternativ inte lagts fram .
Man borde ha betonat att all understödspolitik förkastas och däremot värderas initiativ och ansvar .
Ni framhåller inte åldrandet av befolkningen som kommer att få grundläggande verkningar på vårt samhälles struktur inte bara ur ekonomisk synpunkt utan också på folkhälsoplanet .
Det handlar egentligen om en tyst revolution och i det avseendet väntade jag mig mera i ert meddelande .
Ni betonar slutligen att den europeiska forskningen står i centrum inför vår framtid .
Ni anger emellertid inte vilka medel ni vill sätta in .
De etiska principerna finns också i centrum av denna forskning .
I ert meddelande nämns ingenting .
Herr ordförande , ni vill ge bättre information till medborgarna .
Börja då med att stärka banden med parlamentet : vi är dessa medborgares företrädare .
Fru talman , ärade ledamöter !
Man kan inte annat än instämma i de allmänna linjerna i femårsprogrammet och programmet för år 2000 , som ordförande Prodi har beskrivit med sådan glöd i dag .
I de båda dokumenten betonas starkt behovet av att fastställa nya former för europeisk governance och att i detta syfte omvärdera kommissionens uppgifter med stringentare prioriteringar i strävan mot full sysselsättning .
Detta genom att samordna staternas ekonomiska politik och socialpolitik på ett mer effektivt sätt och - vilket jag tillåter mig att understryka - i första hand de länder som ingår i den monetära unionen och som måste sättas i stånd att utgöra det första exemplet på stärkt samarbete .
I detta syfte nöjer jag mig med att betona tre av de viktiga prioriterade frågor som bör vägleda Europeiska unionens verksamhet under de närmaste månaderna , förutom beträffande kommissionens uppgifter också vad gäller att formulera handlingsprogram för unionens regeringar .
För det första att främja och delta i framtagandet av gemensamma projekt för att skapa ett integrerat servicenätverk inom transport- och energisektorerna , med stöd av Europeiska investeringsbanken .
För det andra att besluta om investeringar som skall genomföras i de enskilda länderna och via gemenskapens projekt inom de prioriterade sektorerna forskning , innovation och uppvärdering av den mänskliga faktorn , som förpliktelser i åtgärdsprogrammen om sysselsättning .
Jag anser att dessa parametrar - särskilt de kvalitativa som är resultat av investeringar i livslångt lärande , fortbildning , anpassningsbarhet och omskolning av de äldsta löntagarna - är mycket mer betydelsefulla och krävande eftersom deras effekter är varaktiga på medellång sikt .
De är något annat än bara uppställandet av årliga kvantitativa mål , som alltid kan ifrågasättas , om att skapa sysselsättning eller minska arbetslösheten .
Om kommissionen bland annat , vilket även understryks i det portugisiska ordförandeskapets program , kunde verka för en ny fas i den sociala dialogen som är inriktad på en överenskommen strategi för social kompetens och kunskapsspridning , kort sagt en strategi för anställbarhet och en definition av reglerna för den , skulle detta göra det möjligt att ta steget till att löntagarna blir informerade och instämmande deltagare i omstrukturerings- och återanställningsprocesserna .
För det tredje tror jag inte att minskningen av antalet aktiva till följd av att befolkningen åldras är ett oundvikligt öde för Europeiska unionen .
Inte bara för att det finns marginaler för att öka kvinnors sysselsättningsgrad och för immigration utan därför att man bestämt måste vända den utbredda tendensen till förtidspensionering och att man tidigt drar sig tillbaka från arbetsmarknaden genom att verkligen inte inrikta den samordnade reformen av de sociala trygghetssystemen på betydande minskningar av de framtida pensionsförmånerna utan på att aktivt utnyttja den ökade förväntade livslängden för att förlänga den yrkesverksamma tiden .
Fru talman , herr kommissionsordförande , mina damer och herrar !
Herr Prodi , ni har trätt in full av ambitioner och reformvilja .
Såväl ni som era ambitioner är välkomna .
De kommer att behövas för den omfattande uppgift vi står inför .
Men för att kunna genomföra alla dessa reformer och driva lagstiftningsprogrammet för år 2001 vidare måste vi vara säkra , inte bara på styrkan hos reformatorn , utan även på de övrigas åsikter .
Ni säger att ni inte kommer att dra er för att komma till oss och be om ökade resurser till kommissionen , men kommissionen bör vara medveten om att vi har en begränsad budget att röra oss med .
Vi förfogar över 1,27 procent av gemenskapens BNI .
Inte en euro mer eller mindre .
Det kommer inte att vara vi som vägrar dessa nya resurser , ni bör då snarare vända er till rådet .
Budgetplanerna är millimeteranpassade .
För att kunna finansiera stabilitetsplanen för Balkanländerna måste man förhandla om den så viktiga granskningen av utgiftsområde 4 , och tänk på de svårigheter vi hade med att godkänna budgeten för år 2000 .
Jag kan påminna er om att vår politiska grupp , PPE-DE , inte tycker om att nya politiska initiativ finansieras på bekostnad av de som redan existerar .
Parlamentet och de europeiska ledamöterna bör fastslå de politiska prioriteringarna .
Tro inte för ett ögonblick att den budgetreform som ni föreslår kommer att dölja begränsningarna av gemenskapens finanssystem .
Det är bra att vi alla i ömsesidigt samförstånd gör en insats för att rationalisera budgeten , men då bör ni vara medveten om att de otillräckliga resurserna , frånvaron av finansiellt självstyre och det bristfälliga genomförandet av budgeten fortsätter att vara angelägna frågor som måste få en lösning .
Därför undrar vi : har kommissionen den politiska viljan att lösa dessa ?
Fru talman , kommissionens meddelande är välskrivet men tillräckligt vagt för att tillåta alla tolkningar .
För det finns ord och därefter deras verkliga politiska betydelse .
Socialdemokraterna applåderar kommissionen när den vill bekämpa social uteslutning och fattigdom .
Men hur skall vi fylla ut gapet mellan politisk retorik och den verkliga världen ?
Vad betyder kommissionens angivna målsättning för en , jag citerar " ekonomisk reform av arbetsmarknaden " ?
Mer flexibilitet , osäkerhet och korttidsanställningar ?
Alla vet att livskvalitet , full sysselsättning och bättre sysselsättning är beroende av en hållbar ekonomisk tillväxt .
Unionen begränsar sig för närvarande till en stabilitetspolitik som förvisso är nödvändig men inte tillräcklig .
Vi socialdemokrater vi önskar få en europeisk pakt för tillväxt och sysselsättning .
Innehållet i denna politik är känt : återupptagande av offentliga och privata investeringar , mer investeringar i forskning , investeringar i grundutbildning och yrkesutbildning och väcka företagsanda .
I det avseendet kan initiativet e-Europa hyllas .
I de nya teknikernas värld är den främsta faran en mer eller mindre lätt tillgång på information beroende på om man är rik eller fattig .
De klyftor som uppstår litet överallt är vår tids främsta problem .
På ena sidan , finns finansmarknadernas överdåd och explosionen av rikedomar medan man på den andra sidan kan notera att uteslutningen ökar .
Man begär att de anställda skall vara flexibla , nydanande och mer och mer produktiva men frukten av denna produktivitet tillfaller mer och mer bara aktieägarna .
Centralbanken är mycket diskret när det gäller finanstillgångarnas överdådiga avkastning men den underlåter aldrig att påminna om att löneökningarna bör vara lägre än produktivitetsökningen .
Hur skall man förklara för de anställda som blir offer för det världsomfattande monopolspelets rationaliseringar att de bör vara beredda att byta yrke flera gånger under sin yrkestid när de stora företagspamparna avgår med ett vederlag på 30 miljoner euro efter att ha förlorat en take-over , som de försökt göra som i poker .
Man har upprepat för oss i åratal att ekonomin måste avregleras .
I de avreglerade sektorerna ser vi nu en mängd fusioner och förvärv som oundvikligen leder till monopolsituationer .
Alla börskamper vilar enbart på i förväg antagna vinstökningar på 15 procent , 20 procent och 25 procent , det vill säga orealistiska procenttal på sikt .
Den tygellösa höjningen av priserna på finansiella och fasta tillgångar betyder att riskerna också ökar .
Den främsta risken som lurar på medellång sikt är inte inflation utan deflation , som kan uppkomma genom att den spekulativa bubblan på de internationella finansmarknaderna spricker .
Fru talman , jag slutar med att säga att de fem kommande åren kommer att vara avgörande .
Det behövs nya regler för globaliseringen , investeringar i realekonomi och i människan .
Staternas synliga hand och kommissionens synliga hand måste säkra marknadsekonomins sociala dimension .
( Applåder ) Fru talman , herr kommissionsordförande , kära kommissionärer , kära kolleger !
Strategidokumentet har enligt min åsikt två tydliga svagheter .
Det hjälper inte att författa en ny ekonomisk och social agenda , när man inte har arbetat av den gamla .
Jag talar om transportpolitiken eller om regionalpolitiken .
För båda områdena har ni med kollegerna Palacio och Barnier utmärkta kommissionärer , och trots detta tillmäter ni dessa områden för liten betydelse i ert strategidokument .
Varför säger jag detta ?
Beträffande transportpolitiken är det viktigt att denna utformas ekonomiskt och miljöpolitiskt förnuftigt i Europeiska unionen , och detta innan andra stater ansluts .
Om kommissionsordföranden lyssnade på mig , så vore jag tacksam , men det är ju inte nödvändigt .
Jag ger er tre exempel på detta .
För det första : Vi behöver en förnuftig avreglering inom järnvägssektorn , ty vi vill föra över godstransporterna från vägarna till järnvägarna .
Det är ekonomiskt och miljöpolitiskt klokt .
Utan avreglering kan vi inte åstadkomma någon förnuftig transportpolitik .
Samma sak gäller den europeiska flygsäkerheten .
Medborgarna har inte någon förståelse för att vi avreglerar lufttransporterna , medan det i luften finns kvar 15 olika sektorer , som kontrolleras nationellt , som medför ekonomiska nackdelar för flyglinjerna och som förstör miljön .
Här måste ni också beta av er föredragningslista .
Herr kommissionär !
Regionalpolitiken nämns alltför litet i ert dokument .
Den sociala och ekonomiska sammanhållningen inom EU är en avgörande uppgift för denna gemenskap .
Om vi inte åstadkommer den , kommer medborgarna i de missgynnade områdena också att vara rädda för utvidgningen .
Vi måste klargöra för dem att vi kommer att använda de närmaste fem åren till att stödja de missgynnade områdena och med en klok användning av medlen göra dem till rika områden .
Då är även de beredda att verkligen rösta för en utvidgning och vara med om att genomföra den .
Herr kommissionsordförande !
Om vi inte lyckas åstadkomma en uttalad solidaritet mellan de rika och fattiga regionerna , då kommer denna union att bli fattigare , och den kommer inte att finna något bifall hos befolkningen !
Herr talman , herr kommissionsordförande , värderade kommissionärer , värderade kolleger !
När vi utformar nya program , får vi inte glömma de äldre program som håller på att genomföras .
Med tanke på detta är det bra att kommissionens arbetsprogram åter tar upp frågorna i Agenda 2000 , den gemensamma jordbrukspolitiken , inklusive fisket , och , för det andra , strukturfondernas verksamhet .
Jag hoppas , herr kommissionsordförande , att detta betyder att den pågående omorganisationen av kommissionen inte kommer att skada den mekanism för kontroll och genomförande som finns i Agenda 2000 .
Frågorna i Agenda 2000 gäller naturligtvis ert tredje och fjärde strategiska mål , den ekonomiska och politiska agendan och den högre livskvalitén .
Vad man kan utläsa av era texter är i vilken utsträckning de högt ställda målen motsvaras av de resurser som kommissionen avser att ställa till förfogande .
Och jag menar inte nödvändigtvis ekonomiska resurser .
För att genomföra Agenda 2000 inom jordbrukssektorn behövs det inte med nödvändighet större ekonomiska resurser , när allt kommer omkring .
Man måste också göra besparingar .
Men det rör sig om intellektuella resurser : man måste investera i humankapital .
Det är nämligen nödvändigt att uppnå två mål , att vidmakthålla den europeiska modellen med ett allsidigt jordbruk , och detta måste ske på ett sätt som underlättar den fria världshandeln med jordbruksprodukter , vilket framför allt gynnar utvecklingsländerna .
Det är inte lätt att kombinera dessa två mål , och det är inte självklart hur det skall gå till .
Eventuellt finns det motsättningar mellan de båda målen , och det finns ingenting som tyder på att kommissionen har uppmärksammat dessa motsättningar och hur de skall lösas .
I fråga om den andra aspekten av agendan , herr kommissionsordförande , den som gäller sammanhållning och regional utveckling , kan vi förvisso uppvisa stora framsteg , men vi har fortfarande efterblivna områden , i synnerhet öområden , som man borde ägna större uppmärksamhet .
Och i fråga om fisket finns det ingenting i ert program som antyder att det rovfiske som hotar att utrota hela fiskarter kommer att få konsekvenser i framtiden .
Det behövs kanske större uppmärksamhet och mera esprit de finesse i dessa frågor .
Fru talman !
Jag vill inleda med att förstärka den varning som många kollegor uttryckt här om denna femårsplan .
När vi lägger fast mycket ambitiösa , långsiktiga mål får vi inte glömma nuet .
Det var något som ledaren för min grupp , Poettering , underströk i sitt inledande anförande .
Unionen skall inte ta på sig en rad nya arbetsuppgifter utan att den centrala grundstommen finns för en framgångsrik europeisk ekonomi .
Den grundstommen är uppenbarligen den inre marknaden .
Hur starkt etablerad är den inre marknaden just nu ?
Jag vill påminna Prodi och de av hans kollegor som fortfarande är här om kommissionens egen undersökning av 3 000 europeiska företag .
Nästan 40 procent av företagen i denna undersökning meddelar att de fortfarande har extra omkostnader för att göra produkter eller tjänster förenliga med nationella specifikationer .
Detta är kommissionens egen undersökning .
Detta är klassiska symtom på att nationella regeringar fortsätter att skapa hinder - byråkratiskt myndighetskrångel som hindrar marknadstillträde .
Kommissionens program visar en störande belåtenhet över genomförandet av den inre marknaden .
Vi måste fortsätta att utöva påtryckningar på alla områden genom att ta bort ytterligare hinder , öka pressen på de medlemsstater som underlåter att sätta den inre marknadens bestämmelser i kraft och naturligtvis utvidga till viktiga nya områden som finansieringstjänster .
Endast med den inre marknaden som stark grundstomme kommer dagordningen för utvidgningen att kunna lyckas .
Ett utvidgat Europa måste byggas på unionens nuvarande starka sidor .
En inre marknad som täcker den utvidgade unionen kommer att vara en fantastisk prestation .
Jag avslutar med att säga på alla mina konservativa kollegors vägnar - och vi är den näst största nationella delegationen i detta parlament - att vi lovar vårt fulla stöd till kommissionen och till Prodi för att de skall lyckas med denna historiska uppgift .
Fru talman , herr ordförande , kära kolleger !
Vid omröstningen om er tillsättning stämde vi möte med er i dag .
Det är nu som de seriösa frågorna börjar , eftersom vi i dag skall uttala oss om ert program .
När det gäller ert inlägg inför kammaren låt mig inrikta mig i mitt uttalande på det som ni kallade det nya ledningssättet .
Ni gör det till ett redskap för försoning med våra medborgare .
Men bakom denna term " nytt ledningssätt " verkar helt enkelt frågan om institutionernas funktion ligga och frågan om våra offentliga myndigheters funktion , om vi är överens om att anse att Europeiska unionen bör vara en offentlig myndighet .
Bandet mellan unionens institutioner , medlemsstaternas befogenheter och de lokala och regionala myndigheterna , det går väl an .
Men är det verkligen så vi kommer att försona medborgarna och den europeiska uppbyggnaden ?
Är det verkligen så vi kommer att svara på de grundläggande frågorna som inte i så hög grad är " vem gör vad " utan snarare " vad gör vi tillsammans " ?
För det är just det som är problemet hos våra medborgare .
I ert uttalande tog ni upp de utmaningar som väntar oss , globaliseringen , utvidgningen och jag vill tillägga framtiden för vår sociala modell .
Därför framhåller vi så starkt med min grupp detta förslag till stadga för det tycks oss att om vi skrev in utformningen av denna stadga om grundläggande rättigheter i vår tidsplan är det just för att vi står vid en historisk mötespunkt , och att unionen behöver omdefiniera de värden kring vilka den byggdes upp inom de aktuella gränserna , men också inför de kommande utvidgningarna som vi önskar så hett , men inte på vilka villkor som helst .
Våra medborgare väntar sig mera Europa av oss , men inte vilket Europa som helst .
De förväntar sig inte att vi skall anpassa oss till globaliseringen , men att vi på grundval av vår sociala modell skall vara en organisationskapacitet för globaliseringen .
Ur den synpunkten bör jag säga er att när ni engagerar er till förmån för en politisk union - och vi är positiva till den politiska unionen - kan detta inte göras om den inte grundas på vår sociala modell och det som utgör vår originalitet och vår kapacitet att bättre styra världens affärer .
Fru talman , herr kommissionsordförande , fru kommissionär , herrar kommissionärer , värderade kolleger !
Jag vill börja med ett citat : " Kommissionen kommer att fortsätta förberedelserna för en europeisk stadga för grundläggande rättigheter och lägga fram förslag för att genomföra ett ambitiöst program .
Kommissionen kommer särskilt att föreslå att en äkta europeisk asyl- och invandringspolitik tas fram , och uttalar sig för att rättshjälpen och rättssamarbetet förstärks och att ett effektivt tillvägagångssätt utvecklas för att bekämpa varje form av brottslighet . "
Detta dokument är en fars i all sin korthet !
En fars därför att vi känner till och uppskattar kommissionär Vitorinos arbete , och det som här läggs fram på papperet står därmed i klar motsatsställning till fakta .
Ett sådant dokument är överhuvud taget inte någon basis för ett poängsystem .
Det har prisats och lovats som en stor prestation , men jag håller fast vid att vi behöver en grund för ett poängsystem .
Vi vill som parlament seriöst diskutera den framtida utvecklingen inom detta politiska område på grundval av ett program .
Det vi förväntar oss är miniminormer i asylförfarandet , för att få snabb hjälp åt flyktingarna men också för att skapa klarhet för dem som inte befinner sig på flykt .
Vi vill ha instrument för att förhindra missbruk .
Vi vill ha en utveckling av invandringspolitiken i gemenskapen , som naturligtvis också inkluderar medlemsstaternas integrationsförmåga , och vi behöver en utbyggnad av exempelvis Europols operativa uppgifter , för att här konkret vidta åtgärder för att bekämpa den organiserade brottsligheten .
Vi befattar oss seriöst och mycket intensivt med dessa uppgifter , och vi förväntar oss samma sak från kommissionens sida , även om de bara handlar om att lägga fram dokument !
Fru talman , herr rådsordförande , ärade kommissionärer , ärade kollegor !
Jag vill ta tillfället i akt och ta upp frågan om Världshandelsorganisationen ( WTO ) , ett område där viss överensstämmelse råder mellan kommissionens dokument och den socialdemokratiska gruppens ståndpunkt , något , som vi redan har hört , inte händer på andra områden .
Det råder en viss överensstämmelse eftersom vi är för ett handelsutbyte på internationell nivå , men vi är för ett sådant handelsutbyte främst tack vare inrättandet av gemensamma lagar , gemensamma regler som kan reglera världshandeln kring ett och samma mål : att handeln skall främja tillväxten , och framför allt att tillväxten blir harmonisk där medborgarnas värde inte bara är något med ensamrätt för de mera dynamiska och konkurrenskraftiga regionerna i världen .
Å andra sidan , vad är det för principer vi vill visa med ett sådant konstaterande ?
På Världshandelsorganisationens nivå har den här regleringen och de här normerna lett till ett ökat handelsutbyte , det vill säga ökad rikedom , men när vi kontrollerar hur rikedomen har fördelats måste vi tyvärr konstatera att avståndet blir allt större mellan världens rikare länder och block och de fattigare och mera underutvecklade länderna .
Därför är vi såväl berättigade som tvungna att ställa oss följande fråga : Vad tjänar de nuvarande gemensamma lagarna till , de nuvarande gemensamma reglerna ?
Vad tjänar de nuvarande förhandlingarna till , såsom de genomförs , och Världshandelsorganisationens nuvarande verksamhet som å ena sidan ökar handelsutbytet , men samtidigt genererar skillnader och ökar avståndet mellan de rika och de fattiga länderna ?
Vi sade därför att vi var positivt inställda till kommissionens strategi inför förhandlingarna i Seattle och följande .
Vi är framför allt för den strategiska visionen , men det krävs mod och djärvhet .
Å ena sidan måste vi kräva att de sociala och miljömässiga rättigheterna samt konsumentskyddet införlivas i de nära förestående förhandlingarna .
Det är dock först och främst fråga om att ha en långsiktig ambitiös och modig vision när det gäller reformen , inte bara av WTO , utan också av Internationella arbetsorganisationen ( ILO ) och Förenta nationerna , men framför allt av de finansiella institutionerna , i första hand Internationella valutafonden ( IMF ) och Världsbanken .
Vi måste vara modiga och inte titta partiskt på globaliseringen , vi måste i stället ha mod att på ett globalt sätt se till att rikedomarna inte bara tillfaller de mera utvecklade länderna , utan alla världens regioner skall få en harmonisk tillväxt och utveckling .
Fru talman !
Även jag vill lovorda kommissionens initiativ att lägga fram en rapport om sina strategiska mål för de närmaste fem åren , även om jag hoppas att man har för avsikt att i senare dokument rätta till det överdrivna antalet generaliseringar och den diffusa prägeln på det dokument som vi behandlar i dag .
Mot bakgrund av detta , fru talman , vill jag än en gång framföra min klagan över frånvaron av en fiskeripolitik .
Det är överraskande att inte kommissionen som ett strategiskt mål för de närmaste åren beslutar om en process med en granskning av denna fråga inom gemenskapspolitiken , inför den reform som bör äga rum år 2002 .
Denna granskningsprocess är , utan tvekan , en av de viktigaste händelser som kommer att påverka fiskesektorn under många år .
Men det verkar den inte vara för kommissionen , som är ansvarig för att innan utgången av år 2001 inför rådet och parlamentet lägga fram en rapport om gemenskapens fiskeripolitik det senaste årtiondet , mot bakgrund av vilken rådet bör fatta lämpliga beslut om en förändring av denna .
Faktum är att en granskningsprocess redan har påbörjats av många yrkesgrupper och institutioner , till exempel av Europaparlamentet , som redan 1998 sammanställde och antog ett betänkande där de aktuella problemen och bristerna inom gemenskapens fiskeripolitik påvisades .
Vi har flera gånger bett om en minimikalender för denna granskning , men vi har inte fått något svar .
Två år minst är ingen lång tid med tanke på den besynnerliga situationen för fiskeripolitiken vad gäller bestämmelserna på den inre marknaden och på att missförhållandena måste lösas inom detta reformförfarande .
Därför ber jag , fru talman , herr kommissionsordförande , att denna fråga , som är av stor betydelse för en så pass viktig sektor inom Europeiska unionen , beaktas i denna strategi och i de strategiska målen för de närmaste fem åren .
Fru talman !
Jag skulle också vilja gratulera till kommissionsordförande Prodis program .
Jag välkomnar särskilt hans erkännande om att denna rättskaffens kammare har upprätthållit tillväxt : informationssamhället på en växande europeisk marknad och dessutom en enda helt fungerande valuta som skall ge oss möjligheten att verkligen främja välfärd , innovationsföretag , entreprenörsandan och - viktigast av allt - arbeten av maximalt varaktigt värde för våra europeiska medborgare .
Jag har en iakttagelse , inte kritik , att redovisa beträffande kommissionsordförande Prodis uttalande i morse som var ganska tandlöst om den ekonomiska politikens verkliga innehåll .
Vi får inte ta någonting för givet i fråga om hur vi kan omstrukturera den europeiska ekonomin .
När allt kommer omkring , vad är social rättvisa om där inte finns full sysselsättning ?
Full sysselsättning är det bästa sättet att skapa social rättvisa för v åra medborgare .
Detta är den centrala fråga som vi skall inrikta oss på .
Jag vill gärna framföra min uppskattning av ett eller två initiativ som kommissionen redan har lagt fram och som skall hjälpa oss : i synnerhet att kommissionär Liikanen förbundit sig att föra en nytänkande kunskapsbaserad ekonomi .
Ja , e-Europa kommer att vara framtiden för oss och hjälpa oss att skapa ny välfärd och nya jobb .
Jag välkomnar kommissionens initiativ nu och tidigare om stöd till våra små och medelstora företag , och jag skulle vilja gratulera vårt portugisiska ordförandeskap för dess initiativ att införa en stadga för småföretag .
Det är viktigt och något som kan behandlas på toppmötet i Lissabon .
Jag välkomnar också kommissionär Busquins idé om att skapa ett gemensamt forskningsområde för hela Europeiska unionen .
Detta är återigen ett sätt för oss att medverka till att skapa bättre möjligheter till sysselsättning och välfärd .
Ni sade i er sammanfattning , kommissionsordförande Prodi , att avreglering , konkurrensmöjligheter , lågt hållen inflation , innovation , vetenskap och teknik är viktiga faktorer för att den europeiska ekonomin skall bli framgångsrik och för att lyckas med att skapa nya jobb i framtiden .
Jag håller verkligen med er om det , men vi kan inte ta något för givet .
Det finns fortfarande mer som vi måste göra och toppmötet i Lissabon skall bli en del av det .
Så med dessa kommentarer vill jag gärna gratulera er till programmet och önska det all framgång .
Fru talman , herr kommissionsordförande !
Jag vill koncentrera mig på två punkter , som inte har nämnts i ert program .
Jag har fått det intrycket att detta strategidokument från kommissionen för de närmaste fem åren skall läsas som ett vetenskapligt arbete om Europeiska unionen , eller som en principförklaring .
Men den ger inte intryck av någon verklig politisk strategi från kommissionens sida .
Som kultur- och utbildningspolitisk talare för min grupp hade jag dessutom av just en italiensk kommissionsordförande kunnat förvänta mig mer innehåll .
På detta vis ger inte kommissionen Europa någon själ !
Det finns inte alls någon kultur eller utbildning i detta dokument .
Men det är nödvändigt att skapa ett verkligt europeiskt utbildnings- och kulturområde .
Bara ett par stickord .
Jag talar om att införliva kulturindustripolitik i detta utbildnings- och kulturområde ; den skapar arbetstillfällen .
Jag talar om att skapa en kulturell mainstreaming på alla politiska områden , om att förstärka och förbättra den europeiska inriktningen på innehållet i utbildningen , liksom om att knyta samman utbildningspolitiken i Europa .
Jag vill understryka det livslånga lärandet .
Herr kommissionsordförande !
Ni talade inte heller om det europeiska audiovisuella området , och detta i början av det nya århundradet !
Dessutom konstaterar jag att informationspolitiken och kommunikationen , som bör anpassas till medborgarnas behov , inte heller nämns .
Jag tror alltså att det fattas något i detta program .
Ett verkligt europeiskt medborgarskap är beroende av att ett verkligt utbildnings- och kulturområde skapas och synliggörs .
Principförklaringar räcker inte !
Vi behöver innehåll som kontinuerligt genomförs av kommissionen på det sätt som jag tidigare förklarade , genom politiska åtgärder .
Fru talman !
Herr Prodi , hur skulle då sammanfattningen av er politik , ert arbetsprogram och er måttstock se ut om ni var tvungen att ställa upp i direkta val ?
Ni har den goda , charmanta idén att resultatet och måttstocken för er politik och för ert femårsprogram kommer att avgöra valresultatet respektive valdeltagandet vid nästa Europaval .
Om jag föreställer mig att jag skall presentera ert arbetsprogram för mina väljare , som jag träffar varje vecka och som jag varje vecka måste förklara det för - inte på högre politisk nivå , utan på gatan - då frågar jag mig vad jag skall säga ?
Herr Prodi , vad skall jag säga att det finns för nyheter i det ?
Det finns ingenting nytt i ert arbetsprogram .
För fem år har ni använt 12 sidor , för ett års arbetsprogram har ni använt 18 sidor .
Ger det mig några förhoppningar för år 2000 ?
Nej , det gör det inte !
I ert arbetsprogram 2000 säger ni något mycket klokt .
Ni säger att miljöhänsyn måste integreras i alla andra politiska områden .
Har ni gjort det , herr Prodi , och har ni också läst årets arbetsprogram ?
Ni har nämligen inte gjort det !
Ni har inte integrerat miljöpolitiken i utvidgningen , fastän det är ett av kärnproblemen i samband med utvidgningen .
Ni har inte heller integrerat den i den ekonomiska politiken , konkurrensen eller den inre marknaden .
Ni har inte gjort det någonstans .
Ni har sammanfogat enskilda sättstycken , men ni har inte skapat någon helhet .
Ni sade tidigare i ert tal att en sådan katastrof som den som skett i Donau måste ge anledning till ett katastrofprogram - nej , herr Prodi , vi måste äntligen börja genomföra lagstiftningen och även se till att vi kan kontrollera lagstiftningen .
Ni skriver i ert femårsprogram att människorna i Europeiska unionen med all rätt förväntar sig bättre livsmedelsstandarder och bättre livsmedelslagstiftning .
Herr Prodi , ni vet inte vad ni talar om !
Europeiska unionens livsmedelslagstiftning är den mest ambitiösa i världen !
Det som saknas , är att den skall genomföras och kontrolleras i medlemsländerna .
Ta äntligen er uppgift på allvar att som ordförande för kommissionen ta medlemsstaterna i öronen och tvinga dem att göra sin plikt och genomföra sina uppgifter !
De skall inte alltid bara ägna sig åt sina fritidssysselsättningar , utan utföra det dagliga normala arbetet .
Det förväntar vi oss av er under de närmaste fem åren !
Fru talman , herr kommissionsordförande , mina damer och herrar !
Ni gör det inte enkelt för mig som ordförande för fiskeriutskottet , herr Prodi .
Jag ser mig tvungen att offentligt här i dag kritisera fiskets frånvaro i det program som ni har lagt fram .
De närmaste fem åren kommer Prodis kommission - detta tillkännager ni högtidligt i den första av era slutsatser - att genomgå stora förändringar .
Jag hoppas att de förändringar som ni tillkännager inte innebär en ännu större diskriminering av fisket , att döma av den väldiga och totala tystnad som frågan omges av i ert program .
Inte en rad , inte ett ord angående fisket eller den gemensamma fiskeripolitiken .
Jag begär inga detaljer eller konkretiseringar , men jag anser att ett omnämnande vore på sin plats .
Hur är det möjligt att en gemensam - jag upprepar , gemensam - politik med en sådan ekonomisk , social och regional genomslagskraft - och som påverkar Europas ekonomiska och sociala sammanhållning , har blivit bortglömd ?
Ännu värre , om möjligt med tanke på att kommissionen , herr Prodi , - så som påpekades - skall genomföra granskningen eller reformen av den aktuella gemensamma fiskeripolitiken , som den är ålagd att göra år 2002 .
Kommer inte kommissionen heller att göra något - åtminstone tillkännages inget sådant - år 2000 åt denna reform ?
Vilket är då budskapet till Europas fiskare , till deras familjer och till fiskeriindustrin , såväl själva fisket som dess bearbetande och saluförande grenar , och till närbesläktade eller stödjande industrier som är beroende av fisket i så och så många europeiska hamnar i så och så många europeiska regioner , många av dem för övrigt i ytterområden , som med all rätt kräver att man fokuserar uppmärksamheten på detta problem ?
Ni hänvisar inför de närmaste åren tydligt till den gemensamma jordbrukspolitiken , men ni säger inget om den gemensamma fiskeripolitiken vad gäller den dubbla anpassning som måste ske av den inre marknaden för att det inte skall finnas några undantag - något som också har påpekats här - i ett globalt sammanhang , i denna globalisering .
Parlamentet har uttalat sig på den första punkten och kommer också att göra det på den andra .
Jag ber er därför , herr Prodi , att ni tar upp detta i ert svar i dag .
Vår parlamentsgrupp kommer att lägga fram ett ändringsförslag i den frågan och jag skulle vilja att ni gav oss ett positivt besked .
Herr kommissionsordförande !
Det här är ett historiskt ögonblick för parlamentet , ett femårsprogram efter kommissionens kris .
Jag skulle för den socialdemokratiska gruppens räkning vilja koncentrera mig på punkten angående inre reformer .
Vi stöder gärna programmet så som det nu lagts fram i en samrådsakt och som även återkommer i vice ordförande Kinnocks program för kommissionens räkning .
Vi tycker det är mycket viktigt att vi , när det gäller ekonomisk kontroll , personalpolitik och kortare byråkrati , ser fram emot snabba beslut och en effektivare byråkrati , till medborgarnas tjänst .
Samtidigt inser vi att det är ett enormt stort program och att under de kommande årens ombyggnad så måste samtidigt butiksförsäljningen fortsätta med konkreta resultat .
På samma sätt som kvinnorna i Nederländerna plötsligt upptäckte att de kunde hänvisa till den europeiska lagstiftningen för att de låg för långt efter med avseende på den sociala tryggheten , gäller i dag också samma sak för flera andra medborgare .
De vill ha resultat .
Demokrati , öppenhet , insyn och tydlighet hör alltid ihop med resultat , medborgare uppskattar resultat och det är på dessa som kommissionen bedöms .
Det är precis som kollega Swoboda och även andra kolleger här redan sagt : rädslan för modernisering , globaliseringen , den enskilda personen som förlorar sin egen trygghet och säkerhet .
Det kan förebyggas med hjälp av den europeiska sociala modellen och om resultat uppnås på alla de här konkreta områdena .
Mitt innerliga yrkande för stöd till den inre reformen hör alltså lika mycket ihop med konkreta resultat på det sociala området , så att medborgaren känner igen sig , här i Europa och även där utanför .
Den medborgaren , en femtedel av världsbefolkningen , har fortfarande inte tillgång till grundläggande sociala möjligheter som till exempel undervisning och hälsovård .
Det är dessa som vi verkligen måste visa solidaritet med .
Fru talman , ärade kommissionsordförande , ärade kollegor !
Jag har läst och återigen läst kommissionens dokument om de strategiska målen för mandatperioden .
Det gläder mig att vi har diskuterat det i parlamentet , jag noterar löftena och jag noterar det som utlämnats .
Kommissionen nämner bara helt apropå den ekonomiska och sociala sammanhållningen , solidariteten mellan medlemsstaterna och Europeiska unionens regionala politik , och detta samtidigt som man tar upp utvidgningsfrågan .
Kan det vara så att målet skall anses vara uppnått med en mindre skillnad mellan tillväxtnivå och det påföljande stödet för den faktiska konvergensen ?
Med all säkerhet inte !
Under tiden menar man mycket riktigt att Europa måste omvärdera rollen som solidarisk partner till u-länderna samt koncentrera sig i kampen mot fattigdomen .
Vad stort sker , det sker tyst .
Kommissionens sätt att inte ta upp sammanhållningen är för mig allvarligt .
Man förringar en princip i fördragen - den ekonomiska och sociala principen - som skall genomsyra all politik och alla åtgärder vidtagna av de europeiska institutionerna , man verkar vara ovetande om att många europeiska regioner är kraftigt underutvecklade , man glömmer att utvidgningen rättfärdigas av ett gott omdöme i den regionala politiken .
Utan verklig konvergens är sammanhållningen inom Europeiska unionen i fara .
Kom ihåg den sjätte periodiska rapporten om tillståndet för Europeiska unionens regioner , som kommissionen är ansvarig för .
Med en genomsnittlig tillväxtnivå på 100 konstaterar man att de tio regioner som anses vara de " starkaste " i genomsnitt ligger på 158 , och de tio " svagaste " stannar på 50 .
Dra era egna slutsatser .
50 : just den tillväxtnivå som min region , Azorerna , hamnade på - en av dem som i fördragen definieras som en ultraperifer region .
Jag väntar på kommissionens betänkande om ultraperifera regioner som rådet fastslog skulle utarbetas till december 1999 .
Jag slutar med att på nytt påtala min övertygelse : utan ekonomisk och social sammanhållning kommer ingen sammanhållning alls att uppnås , bara upplösning .
Fru talman , herr ordförande !
Vi och den europeiska allmänheten behöver en stark kommission , för enligt fördragen och också folkets vilja är kommissionen motorn i den europeiska uppbyggnaden , den Sisyfosklippa som vi tillsammans måste bära upp till toppen igen efter varje utvidgning .
Således , en stark kommission men som stöder sig på parlamentet , och parlamentet är således er allierade , men det är en besvärlig allierad vars meddelanden bör avlyssnas och jag skulle vilja lämna några meddelanden i detta korta inlägg .
För det första , herr ordförande tror jag att även om era båda föregångare huvudsakligen ägnade sig åt att utveckla en inre marknad och inrätta en gemensam valuta är det huvudsakligen er sak att utveckla det medborgarvärde som står i centrum för den europeiska uppbyggnaden .
Ni får nämligen inte låta er distraheras enbart av utvidgningsärendet , hur viktigt det än är .
Ni måste gå längre i riktning mot en försoning av medborgarna med Europa och i synnerhet de medborgare som är offer för ekonomiska , sociala och otvivelaktigt på sikt tekniska brytningar .
Främjandet av vetenskaplig utveckling , även främjandet av nya tekniker och allas tillgång till dessa tekniker kommer inte att säkras av marknaden och av konkurrensen , inte mer än att marknaden och konkurrensen kommer att säkra den sociala närheten och effektiviteten när det gäller de stora kollektiva tjänsterna , hälsa , utbildning , transporter , kommunikationer , vatten och jag vet inte vad .
Ert åtgärdsprogram och era målsättningar är diskreta och rentav helt tysta när det gäller konsolideringen och finansieringen av de stora offentliga tjänsterna och tjänster av allmänt intresse .
Det finns en absolut prioritering , herr ordförande , om ni vill försona Europa med medborgarna : att se till att de hellre väljer Europa än Jörg Haider .
Fru talman !
Kommissionen gjorde rätt när den gjorde livsmedelssäkerhet till en av de viktigaste frågorna .
Den nyligen inträffade dioxinskräckhistorien i Belgien , den tidigare BSE-krisen i Storbritannien och den pågående kontroversen om hur farliga genetiskt modifierade livsmedel är har alla bidragit till att konsumenterna litar mindre på att den mat de äter är ofarlig .
Om kommissionen verkligen kan återställa förtroendet för livsmedelsproduktionskedjan kommer den samtidigt att återskapa förtroendet för Europeiska unionens institutioner och visa deras förmåga att skydda EU-medborgarnas rättigheter .
Jag välkomnar därför det faktum att frågan om livsmedelssäkerhet , folkhälsa och konsumentförtroende understryks markant i kommissionens arbetsprogram för år 2000 .
Jag blev dock besviken över hur förslaget om inrättandet av en europeisk livsmedelsmyndighet är utformad i den senaste vitboken .
I dess nuvarande form är det som föreslås mer som ett rådgivande organ till kommissionen snarare än ett självständigt organ som skulle ha beslutande och lagstiftande befogenheter mer likt dem hos den amerikanska livsmedelsmyndigheten : Food and Drug Administration , vilken redan har skapat trovärdighet på detta speciella område .
Vidare måste man i det framtida lagstiftningsarbetet ta itu med arbetsmetoden för samspelet mellan den europeiska livsmedelsmyndigheten och myndigheterna i nationella medlemsstater , exempelvis myndigheten för livsmedelskontroll i Irland .
Detta organ , exempelvis , utför tillsammans med det nyligen inrättade gränskontrollorganet i Irland för livsmedelssäkerhet redan ett bra arbete .
Det skulle vara tragiskt om deras ansträngningar skulle undergrävas på grund av brister i EU : s lagstiftning .
Jag fruktar att sådana brister i EU : s lagstiftning kan leda till revirstrider mellan nationella organ och EU-organ , som borde arbeta tillsammans i stället för att mot varandra .
Det är något som vi måste bevaka .
Fru talman !
Ordförande Prodis presentation i dag var nödvändigtvis en ganska brett svepande historia .
Vi kommer att titta efter enskilda detaljer år för år , till exempel i det sociala åtgärdsprogrammet som skall läggas fram i år .
Vi skall också granska detta från perspektivet social- och sysselsättningspolitik och genomföra en rad kontroller .
Vi skall granska i vilken omfattning vi kan skapa en liksidig triangelformad politik där man kombinerar ekonomisk politik , sysselsättningspolitik och socialpolitik .
För ögonblicket ligger socialpolitiken långt bakom politikområdena ekonomi och sysselsättning .
Inom ramen för sysselsättningsstrategin skall vi sträva efter att fördjupa och bredda strategin efter översynen under det portugisiska ordförandeskapet och inom den ram som förslagits av det portugisiska ordförandeskapet .
Inom ramen för den sociala dimensionen skall vi sträva efter att fördjupa den inre marknaden med en social aspekt .
Strömmen av sammanslagningar , fusioner och överlåtelser som vi upplever när marknaden får allt större intresse innebär att vi måste göra något för att aktualisera den mall för de informations- och samrådsdirektiv som vi antagit tidigare ; men vi måste också komplettera dem med det nya generella regelverket för information och samråd och uppdatera företagsrådsdirektivet .
Vi behöver även en uppförandekod för bolag för att se till att företag i själva verket arbetar i partnerskap med sina anställda i förändringsarbetet .
Det är ett framgångsrikt sätt att hantera förändring och jag hoppas kommissionen kommer att se till att det genomförs .
Slutligen , med uppdykandet och återuppvaknandet av rätten till främlingsfientlighet inom Europeiska unionen hoppas jag att våra institutioner tillsammans kommer att göra sitt yttersta för att ge artikel 6 verkligt innehåll genom att tillämpa artikel 13 för att bekämpa diskriminering och artikel 137 för att bekämpa uteslutning .
Vi måste snarast börja arbeta med den dagordningen nu .
Förhoppningarna , ordförande Prodi , är bra men vi vill att dessa förhoppningar skall paras med åtgärder .
Fru talman !
Jag hoppas att det är ett gott tecken att jag avslutningsvis får påpeka ytterligare en sak !
Herr Prodi , i era reformsträvanden är ni särskilt intresserad av att förverkliga en framtidsorienterad sysselsättningspolitik över hela Europa .
Men för just den ekonomiska sektor som jag företräder , fiskerisektorn , betyder detta förändringar .
Vi måste överge de planekonomiska subventionerna och komma fram till en liberal politik , som främjar det egna ansvaret .
Vi måste sänka skyddstullarna för att garantera att företagen inom tillverkningsindustrin tas i anspråk effektivt .
Så handlar det slutligen om det europeiska näringslivets konkurrenskraft på världsmarknaden och om tusentals arbetstillfällen inom tillverkningsindustri och havsfiske .
Men jag behöver säkert inte påminna er om betydelsen av en näringsgren som inte bara är en nationalekonomisk faktor , utan också en samhällsfaktor , som inte bara berör Tyskland , utan gränsövergripande berör alla kustregioner i Europa .
Dessutom är denna näringsgren en av de få sektorer som fullt ut har integrerat europeiskt besluts- och handlingsansvar .
Därför förväntar vi också här att vi får medbeslutanderätt .
Det rekommenderas nu enhälligt .
Men revideringen av fiskeripolitiken är fastställd till att äga rum om några månader , dvs. i början av år 2000 .
Då är det verkligen störande att denna näringsgren alls inte nämns i föreliggande dokument .
Jag hoppas att det här handlar om ett missförstånd !
Jag ber , herr Prodi , att stå för vad ni sagt , och genomföra det !
Fru talman !
Många av talarna från socialistgruppen har redan identifierat viktiga områden där det finns brister i kommissionens uttalande .
Vi har dock uttryckt att detta är ett nyskapande och mycket välkommet initiativ av kommissionen .
Ett område som jag vill inrikta mig på , förutom dem som redan nämnts , är kulturell mångfald i Europa .
I inledningen till detta uttalande tillstås i avsnittet om livskvalitet att detta är viktigt .
Men det finns inget i uttalandet som visar att kommissionen avser att vidta några åtgärder för att hantera frågan om kulturell mångfald .
Om vi skall kunna garantera att vi besegrar dem som sprider rädsla ibland oss - dem som strävar efter makt med stöd av oroliga medborgare - då måste vi allvarligt ta itu med frågan om hur vi kan leva tillsammans och hur vi kan undanröja de negativa stereotyper som vi har om varandra , både inom den nuvarande Europeiska unionen och bland dem som försöker ansluta sig och rent av bland dem i andra delar av Europa och världen som vill komma hit och bo och arbeta i Europa .
Om vi inte tar itu med dessa frågor , om vi inte kan undanröja dessa negativa stereotypa uppfattningar , om vi inte använder det som är bäst från våra olika kulturer och språk och skyddar och utökar det och ser till att vi menar allvar med att ha ett mångfaldigt Europa , kommer vi att misslyckas .
De som just nu är i blickpunkten i Europa grundat på rädsla skall vinna slaget .
Jag är allvarligt oroad att om kommissionen inte inser att detta är en viktig aspekt på hur vi skall skapa ett samhörande Europa kommer vi att göra framsteg på det ekonomiska området och på sysselsättningsområdet och även inom utrikes- och säkerhetspolitik men våra medborgare kommer fortfarande att vara ängsliga därför att de kommer att vara rädda för det okända och rädda för dem som de inte förstår .
Om vi inte vidtar åtgärder för att hantera detta kommer vi till sist att misslyckas .
Kära kollega , jag tackar er .
Innan jag på nytt ger ordet till kommissionens ordförande vill jag meddela er att jag i enlighet med artikel 37 har fått sju resolutionsförslag till sammanfattning av debatten . .
( IT ) Fru talman , ledamöter !
Jag tackar er för denna kraftfulla , seriösa och konstruktiva debatt .
Det har varit en fredlig debatt med en stor samsyn om de grundläggande punkterna , men även med en bred bekräftelse av parlamentets rättigheter och behovet av samarbete och konfrontation mellan parlamentet , kommissionen och rådet .
Det har varit en konstruktiv debatt för vårt Europa .
Det har sagts att det dokument vi har framlagt är ett politiskt manifest som innehåller vissa inre motsägelser .
Fru Hautala , jag tror nästan att ni som sade detta har rätt , för mitt dokument är faktiskt ett politiskt manifest .
Men det är inget abstrakt politiskt manifest , det är ett manifest om en politisk vilja som vi behöver i denna känsliga fas för Europa .
Det tjänar ingenting till att säga att Europa är i kris om vi sedan inte klarar av att lägga fram ett politiskt manifest , diskutera det , slåss om det och gå vidare tillsammans med slutsatserna av detta .
De motsägelser som sedan Hautala rätteligen har noterat mellan mål och medel är de motsägelser som finns i den aktuella europeiska verkligheten , de motsägelser som vi är kallade att sanera och komma över : detta är vidden av den politiska uppgift vi har i dag .
Jag har belyst dessa motsägelser utan att dölja något : det gläder mig att de har betonats så väl och även ibland framhävs maximalt och det är därför vi vill förändra de instrument som styr vår verksamhet , parlamentets verksamhet , min verksamhet , alla de europeiska institutionernas verksamhet .
Det är därför vi ville ha en stark regeringskonferens och därför som Helsingfors var en känslig fas .
Man har skrivit att vi har låtit bli att driva på för ett starkare Europa och sedan har det visat sig att vi tvärtom i Helsingfors lyckades hålla en låga brinnande som sedan har tagit sig ännu mer .
Tänk på det tal Republiken Frankrikes president höll - jag hänvisar till det här för att det hölls i just denna kammare - om problemen med ett utökat samarbete som återupptog en dialog som tidigare verkade avslutad .
Jag hoppas att den ihärdighet med vilken vi har hållit fast vid ståndpunkterna från Helsingfors kommer att få sin belöning under regeringskonferensen som skall avslutas vid toppmötet i Nice .
Alla - inte bara ledamöterna Poettering och Fiori , utan många talare - har hänvisat till globaliseringen och de svårigheter den medför för våra liv och vår politik .
Kommissionen vill ha globaliseringen , anser att den är positiv eftersom den för upp miljarder människor som var utslagna från världsmarknaden på en miniminivå av anständighet .
Det är tack vare denna globalisering som Kina och Indien och , jag upprepar det , några miljarder människor håller på att vakna .
Jag hoppas att globaliseringen även i framtiden kommer att ha detta positiva innehåll , men den skapar problem i de fattiga länderna och i våra länder , problem vi måste ta itu med .
Detta kommer att bli en av våra stora uppgifter i framtiden .
Den skapar också problem inom de svagaste kategorierna i våra länder .
Det är en rannsakning av våra samveten som vi , dag för dag , måste göra om de verksamma faktorerna , eftersom det står klart att globaliseringen skapar klyftor i våra samhällen , ökar vår fattigdom , ökar mycken ilska , orsakar indelning och uppdelning inom lönenivåer , även för kategorier som verkade homogena , och på detta måste vi fokusera vår uppmärksamhet .
Det är klart att våra unga nyutbildade akademiker konstaterar att det finns löneskillnader som är mer eller mindre stora beroende på den anställning de får och när finanssektorn erbjuder löner som är x gånger högre än för den som till exempel arbetar med forskning , skapar detta problem för hur vårt framtida samhälle skall organiseras .
Detta måste vi fundera ingående över och ärligt talat - och med detta svarar jag Trentin - har vi inte ännu , åtminstone har inte jag ännu , förberett ett heltäckande svar på detta .
Jag började svara i Lissabon , och försökte minska utslagningen av en hel åldersgrupp genom att ombesörja nya kommunikationsredskap för alla unga i Europa , förena alla Europas skolor under en flagg , skapa nya möjligheter för att förhindra geografisk utslagning och utslagning av samhällsgrupper i Europa .
Det är fortfarande för litet för att kontrollera globaliseringen , eller åtminstone förstå dess konsekvenser , men det är ett kraftfullt svar och ett svar vi måste ge .
Det finns också ett svar på global nivå som kommissionen med kraft har framfört under de senaste veckorna via kommissionär Lamy : att återställa förtroendet för tillväxt i tredje världen , som så allvarligt sattes på spel i Seattle , att återskapa WTO : s roll med en omfattande dagordning som just kan klara utmaningen från globaliseringen .
Kommissionen föreslog i Geneve ett kortsiktigt paket som är ovanligt modigt och går många av era krav till mötes .
Vi föreslog ett ensidigt slopande av tullarna för de 38-40 fattigaste länderna , unilateralt , totalt , generellt .
Vi föreslog en reformering av WTO : s rutiner och ökad insyn och vi föreslog att man svarar utvecklingsländerna om problemen med att utöka denna åtgärd .
Om dessa åtgärder kommer vidare under de närmaste dagarna kommer kommissionen - som vi redan har flaggat för - att med kraft driva en nylansering av rundan i sommar , alltså en ny omgång .
Vi försöker sy ihop det sår som öppnades i Seattle .
Detta är kommissionens stora uppgift och samtidigt ett förslag till reformering av WTO med kommissionens bistånd där man äntligen analyserar frågan på djupet , för det har aldrig gjorts under dessa år .
Detta är ett första konkret svar i ett femårsprogram , som inte är till för att ge svar i enskilda frågor utan för att ge just dessa stora linjer , dessa utdrag ur vår framtida verksamhet , utdrag där parlamentets kontroll är viktig och där samarbetet mellan parlamentet och kommissionen är viktigt .
Synergieffekterna mellan kommissionen , parlamentet och rådet är avsevärda , ledamot Cox .
Det står klart att detta tvingar oss att omvärdera konceptet subsidiaritet , som vi har sett och vilket en stor del av mitt inlägg handlade om .
Jag är tacksam mot ledamöterna Poettering , Cox och de andra som har tagit upp det .
Detta är programmets hörnpelare .
Subsidiariteten har alltför ofta betygats vördnad i abstrakt mening men inte tillämpats konkret .
Vi måste ge subsidiariteten ett konkret ansikte och en politisk själ : detta är syftet med vitboken , som skall återge Europa dess värde och ange de konkreta åtgärder som skall genomföras .
Jag vill inte sälja ut Europa , ledamot Dell ' Alba , jag vill inte nedrusta genomförandet av den gemensamma politiken .
Tvärtom vill jag förstärka , påskynda och förbättra besluten och genomförandet av den gemensamma politiken , men jag vill samtidigt undvika att våra system skär ihop på grund av ett stort antal politiska fragment som egentligen inte har mycket gemensamt .
Låt oss komma ihåg hur många gånger vi har gjorts till åtlöje för att vi ägnar oss åt saker som är fullständigt löjliga , som motsäger det sunda förnuftet och motverkar vår befolknings intressen .
Kommissionen kan och måste verkligen vara en föregångare på detta område och för denna omvandling och avlastas onödiga bördor och bli mer trovärdig eftersom den ägnar sig åt core business , eftersom den inte begär utan vägrar ta på sig onödiga uppgifter och befogenheter .
Kommissionen måste bli en pådrivande kraft .
Som Cox sade , " enabling Europe " och inte " including Europe " , och många gånger har vi varit å ena sidan enabling och å den andra including .
Försäkran nummer två : dessa är inte tomma föresatser .
Vi har redan börjat arbeta på dem , inte bara för den interna reformeringen av kommissionen tillsammans med kommissionär Kinnock , utan även i några första reformer av politiska sakfrågors uppbyggnad .
Vi skall ge er ett exempel : om det finns något politiskt område som ligger kommissionen varmt om hjärtat så är det konkurrenspolitiken .
Nåväl , vi har lagt fram ett förslag till reform - och denna kammare stödde denna idé med mycket stor majoritet i januari - som skall möjliggöra för kommissionen att koncentrera sig på kampen mot de allvarligaste konkurrensbrotten , de som är mest framträdande på europeisk nivå , och inom detta område har vi startat ett bredare samarbete än de nationella myndigheterna .
Detsamma har vi gjort om vitboken om livsmedel .
Jag har hört kritik - och jag förstår kritiken - om att " den har mindre makt än den amerikanska Food and Drug Administration " .
Ja visst !
Jag ville utnyttja de nationella myndigheterna som redan är verksamma på området .
Om jag skulle ha använt ett organisationsschema som det amerikanska hade ni gjort uppror i dag och sagt : " Ni har skapat ännu en centraliserad maktapparat i Bryssel ! "
Detta är Europa : denna ömtåliga jämvikt mellan de nationella strukturer som finns i dag och som måste värdesättas , sättas in i ett nätverk med den europeiska myndigheten , inte förödmjukas av att en europeisk myndighet tillkommer .
Det är en svår utmaning eftersom man hittills aldrig har försökt sig på det , liksom utmaningen med utvidgningen är svår .
Jag uppskattar den stora enigheten om utvidgningen .
Det har knappt hörts en enda skiljaktig mening i debatten i förmiddag , och jag uppskattar det eftersom utvidgningen kommer att bli ett beslut som medför uppoffringar för oss , som medför stora förändringar hos oss själva .
Vid tidpunkten för det konkreta beslutet här måste vi och ni stå eniga för att visa att utvidgningen ligger i fredens och välståndets intresse och genomförs som en garanti för våra folk , liksom för de länder som försöker utvidga sig , som jag sade tidigare .
Jag har inte en tanke på att gå vidare med en utvidgning som inte är seriös , som inte är stark , och framför allt - ledamot Muscardini var mycket uppmärksam och gjorde ett riktigt påpekande - kan inte utvidgningen skapa två sorters medlemmar : Utvidgningens förnämlighet ligger just i det faktum att när ett land väl kommer in här är det jämställt med alla de andra .
Jag sade att vi är ett förbund av minoriteter , en union av minoriteter : detta är det fantastiska med Europeiska unionen .
Men utvidgningen består också av stränghet .
Man har påmint mig om problemet med kärnkraftverken och problemet Donau .
De senaste dagarna har jag varit i Litauen , Slovakien och Rumänien : tre länder där vi har tvingats begära att kärnkraftverk skall stängas .
Det har vi gjort medvetna om de allvarliga problemen för de lokala ekonomierna , men vi har förklarat att detta är Europas regler , vi har förklarat att det är en säkerhetsåtgärd som alla bör vidta , som alla måste vidta , som alla vidtar .
Detta har dessa länder som vi har hjälpt med omställningen förstått .
De har engagerat sig i stängningen av kärnkraftverk , som är en enorm uppoffring för dem .
Men detta är Europa : Varför uppoffra sig ?
För att det mål som ligger i allas gemensamma intresse skall uppnås .
Jag tror att det är viktigt att vi finner en samsyn även om Afrika .
Jag har hört många brinnande inlägg om Afrika , som även jag tog upp i mitt anförande för Afrika är ett kors för oss : ingen bryr sig om Afrika .
Jag påminner om den stora rundresa den amerikanske presidenten har gjort under de senaste åren , som gav en strimma av hopp , sedan följde ingenting av detta .
Afrika är i huvudsak vårt problem .
Det finns naturligtvis med i den utrikespolitiska analys vi gjorde förut : frågan om utvidgning , Medelhavet , Ukraina , Ryssland och detta afrikanska problem som vi tittar på .
Förberedelserna för toppmötet går framåt , men det finns enorma svårigheter : det finns dramatiska skiljelinjer i Afrika , och jag försöker även i denna mening minska dem , jag försöker laga sprickor som en nödvändig förutsättning för att skapa en stor politik för detta så desperata Afrika .
Task force vid GD Bistånd arbetar i nära samarbete med GD Yttre förbindelser för att också verka inom nya områden i Afrika .
Vi börjar samarbeta inom kommunikationer , utbildning och vetenskap .
Om vi inte sätter fart inom dessa civilisationsområden kan inte Afrika göra det .
Jag är dock medveten om att vi fortfarande befinner oss i början och ber därför om stor öppenhet och stor hjälp med detta .
Man har också förebrått mig för att jag inte tog upp vissa viktiga kapitel som fisket .
Det är riktigt , jag tog inte upp fisket .
Jag tog inte heller upp jordbruket eller skolan och jag tog inte upp hela den stora äldrevårdspolitiken .
Jag tog inte upp det eftersom jag tycker att en femårsplan skall ge de stora riktlinjerna för utvecklingen generellt sett , men jag är övertygad om dess enorma vikt för den europeiska sammanhållningen och solidariteten .
Jag försäkrar er om ett engagemang på detta område eftersom det är klart att det ingår i läggandet av den storslagna mosaik vi har skisserat i debatten i dag .
Kommissionen måste lägga manken till , just inom dessa våra huvudfunktioner där vi måste göra vår oersättliga roll som politisk och moralisk ledare för Europa gällande för att visa på fördelar och kostnader med vår politik , för att vara mycket tydliga gentemot befolkningen som kräver tydlighet av oss , som kräver total insyn .
På denna punkt lugnar och uppmuntrar mig denna debatt .
Den lugnar mig eftersom jag har uppfattat en bred samsyn om de grundläggande dragen i vårt program , och eftersom jag har intrycket att man har förstått dess verkliga innehåll .
Det har varit en fredlig debatt , som jag sade i början , men inte avslagen , tvärtom har det varit en debatt med enbart hög politisk profil .
Så om termen " manifest " kan ha en negativ klang , äger den dock också stor giltighet , ett starkt politiskt innehåll .
Vi har talat med ett språk som Barón Crespo kallade rakt och öppet .
Det har framkommit klart , men med kraft , att vad vi har framför oss är de stora politiska utmaningar vi måste ta itu med tillsammans .
Detta gör ett intimt samarbete mellan parlamentet och kommissionen än viktigare .
Det får mig att känna mig uppmuntrad .
Somliga blev inte övertygade av anförandet , som Wurtz som i sitt uttalande sade att han uppskattade den konstruktiva andan och som också sade : " Vi har fem år på oss att lyckas " .
Vi är beredda att samarbeta .
Det är det jag vill , och inte - Cox - för att jag någonsin har märkt att jag upplevde en smekmånad .
Ni sade att smekmånaden är slut .
Mina minnen från min smekmånad är något annorlunda än från de månader vi har tillbringat tillsammans , men det gläder mig att ni använde detta ord .
Hur som helst går jag ur denna debatt än mer övertygad om att de stora utmaningar som väntar oss är politiska utmaningar .
De fordrar stor energi , en energi som kommer att bli större ju större synergieffekterna mellan institutionerna blir .
Jag skulle vilja avsluta med den hänvisning Barón Crespo gjorde .
Han hänvisade till någonting som är mig mycket kärt när han nämnde Ambrogio Lorenzettis fresk om det goda styret i Siena .
Om ni minns den är det är en fresk där allting fungerar .
Det finns människor som arbetar , det finns handel , det finns hierarkier som man känner igen mycket klart i samhället Siena .
Det var en veritabel femårsplan för Sienas kommun .
Det var deras dokument med vilket de ville spegla samhället som det var .
Vi kan inte känna annat än beundran , för egentligen kan den vara en riktpunkt .
Ledamot Barón Crespo , vi får inte heller glömma bort att femårsplanen inte kan ha haft något inflytande på världen i praktiken .
Den försvann från de politiska manifesten när Sienas roll i världen försvagades .
Jag tror att vi bör undvika denna fara .
( Applåder )
 
Välkomsthälsning Jag vill meddela att en delegation från Kuwait , som leds av Hans Höghet shejk Salem Al-Sabah , vice premiärminister och försvarsminister är närvarande på hedersläktaren .
På Europaparlamentets vägnar önskar jag er välkomna .
( Applåder ) Herr talman !
Jag skulle vilja ta upp en ordningspunkt som gäller de aktiviteter som i dag organiserades av föreningen för parlamentariska assistenter för att få stöd för sitt krav om att en stadga för assistenter antas så snart som möjligt .
Jag har uppfattat att den 26 januari skrev föreningen till kvestorskollegiet och begärde tillstånd att ställa upp ett bord utanför kammaren i dag för att presentera sitt initiativ .
Samma dag , har jag förstått , gav Balfe assistenterna tillstånd att göra detta .
Sessionstjänsten bad att få träffa assistenterna i går för att gå igenom de praktiska arrangemangen .
Mötet inställdes dock i sista minuten .
Parlamentet har ännu inte meddelat varför tillståndet drogs tillbaka .
Banotti lovade uppenbarligen att skriva ett brev och förklara varför tillståndet drogs tillbaka men hittills har man inte mottagit något brev .
Kan ni förklara varför det tillstånd som gavs till assistenterna drogs tillbaka i sista minuten ?
Håller ni med om att assistenterna driver ett legitimt ärende som måste få höras ?
Kommer ni att göra allt ni kan för att se till att sådant inte kan hända på nytt ?
Kommer ni att göra allt ni kan för att se till att en stadga för assistenterna antas så snart som möjligt ?
Slutligen kommer ni under tiden se till att parlamentets bestämmelser verkligen iakttas och att assistenterna får betalt , som de borde bli , på basis av allt det arbete som de gör för oss ?
Utan dem skulle vi inte kunna sköta våra arbetsuppgifter .
( Applåder ) Herr talman !
Även jag vill ta upp en ordningsfråga .
Finns det några regler eller förordningar som reglerar demonstrationer inom parlamentets byggnad , utanför dörrarna till kammaren , för att säkerställa att ledamöter kan komma in i denna kammare för att fullgöra sina uppdrag ?
Om det finns sådana regler vem ansvarar för att de efterlevs och vad gör de för att uppfylla det ansvaret ?
Herr talman !
Jag skulle vilja ta upp frågan om assistentstadga igen , som vi alltid har prioriterat , och informera er om att vi - den italienska delegationen i gruppen - på gruppens ordförande Barón Crespos uppmaning har deponerat de kontrakt vi har upprättat med assistenterna hos kvestorerna .
Jag tycker att det är en konkret gest för att komma till en lösning på detta problem .
Därför skulle jag vilja uppmana parlamentets presidium att överväga om det inte vore lämpligt att presidiet uppmanade alla ledamöterna att göra detsamma .
Herr talman !
Låt mig först och främst säga att jag helt stöder kravet på en stadga för assistenter .
I går när jag anlände till parlamentet fick jag en skrivelse om en föreslagen demonstration av assistenterna utanför parlamentets dörrar .
Som alla kollegor känner till - och många av er har kontaktat mig under de senaste sex månaderna - bedöms alla utställningar och liknande arrangemang först av parlamentets Comartkommitté ( Comité des Arts - konstkommittén ) .
För att ge ett ej omtvistat exempel : inga kommersiella utställningar får hållas här i parlamentet av uppenbara skäl .
Efter att jag mottog ett brev i går informerade jag omedelbart assistenterna att vi skulle föreslå att de fick hålla ett möte eller demonstration , förmodligen inom en snar framtid och eventuellt under nästa månad .
Men alla sådana arrangemang måste genomföras på ett sätt som inte stör parlamentets reguljära verksamhet .
Jag undertecknade ett brev i går eftermiddag vid parlamentspresidiets sammanträde i vilket assistenterna informerades om detta .
Men jag har också hört att de informerades muntligen om detta beslut av gruppordförandekommittén i torsdag , så de var helt medvetna om beslutet .
Problemet är inte att de talar om för oss hur de känner , det är inga problem med ett eventuellt möte under parlamentets nästa delsession .
Men det blev ett missförstånd då de mottog ett brev från en annan person som de ansåg gav dem tillstånd .
Alla utställningar blir emellertid först bedömda av den så kallade Comartkommittén .
Som ni vet har vi många utställningar runt om i parlamentsbyggnaden om olika länder eller om vad som helst .
Detta är inte ett försök att vare sig censurera eller gå emot den mycket reella och befogade principen att vi bör ha en stadga för assistenter .
Tack för det , ledamot Banotti .
Ert inlägg borde kunna klargöra olika frågor som har tagits upp .
Herr talman !
Jag vill understryka en viktig principfråga .
Personligen anser jag att det är inget mindre än skandal att vi har ledamöter i detta parlament som angriper demonstrationen hellre än att söka lösningen på problemet , vilket är rimliga arbetsförhållanden , rimlig lön och rimliga arbetstider .
( Vi skall nu genomföra omröstningen.1
 
OMRÖSTNING ( Förfarande utan betänkande ) ( Parlamentet godkände förslaget . )
Resolutionsförslag ( B5-0095 / 2000 ) " Området med frihet , säkerhet och rättvisa " ( Parlamentet förkastade resolutionsförslaget . )
Resolutionsförslag ( B5-0109 / 2000 ) " Området med frihet , säkerhet och rättvisa " ( Parlamentet godkände resolutionen . )
Betänkande ( A5-0026 / 2000 ) av McCarthy för utskottet för regionalpolitik , transport och turism om meddelandet från kommissionens till medlemsstaterna om fastställande av riktlinjer för ett gemenskapsinitiativ för ekonomisk och social förnyelse av städer och förorter som befinner sig på tillbakagång för att främja hållbar stadsutveckling ( Urban ) ( KOM ( 1999 ) 477 - C5-0242 / 1999 - 1999 / 2177 ( COS ) ) ( Parlamentet godkände resolutionen . )
Betänkande ( A5-0028 / 2000 ) av Decourrière för utskottet för regionalpolitik , transport och turism om kommissionens meddelande till medlemsstaterna med riktlinjer för ett gemenskapsinitiativ som rör transeuropeiskt samarbete som syftar till en harmonisk och balanserad utveckling i Europa ( Interreg ) ( KOM ( 1999 ) 479 - C5-0243 / 1999 - 1999 / 2178 ( COS ) ) ( Parlamentet godkände resolutionen . )
Betänkande ( A5-0024 / 2000 ) av Procacci för utskottet för jordbruk och landsbygdens utveckling om förslaget till kommissionens meddelande till medlemsstaterna om fastställande av riktlinjer för gemenskapsinitiativet för landsbygdens utveckling ( Leader + ) ( KOM ( 1999 ) 475 - C5-0259 / 1999 - 1999 / 2185 ( COS ) ) 1 .
Röstförklaringar Resolutionen " Området med frihet , säkerhet och rättvisa " Berthu ( UEN ) .
( FR ) Den resolution som parlamentet just har godkänt trots de negativa rösterna från Gruppen Unionen för nationernas Europa om invandringspolitiken styrker retroaktivt den fruktan som vi uttryckte vid ratificeringen av Amsterdamfördraget .
Europaparlamentet visar i fråga om innehållet den mest totala släpphänthet och begär på samma gång mer och mer beslutandemakt till nackdel för de nationella parlamenten .
Sammantaget utgör dessa båda ståndpunkter en blandning som skulle kunna bli katastrofal för Europa på sikt .
När det gäller innehållet har jag i resolutionen räknat till inte mindre än sju uppmaningar på olika ställen om lika rättigheter mellan medborgare i länderna i Europa och lagliga invandrare .
Det är en riktig plåga .
Vad beträffar kampen mot olaglig invandring intresserar det knappast parlamentet .
Det sägs absolut ingenting i resolutionen om gränskontroll och när frågan om Eurodac eller avtalen om återtagande berörs helt kort är det för att beklaga rådets alltför stora fasthet i dessa avseenden .
Däremot saknas inte den traditionella maningen att bilda en fond för flyktingar som skall finansieras med gemenskapens budget .
Europaparlamentet begär slutligen att invandringspolitiken skall ses över i förhållande till den demografiska situationen .
Man vet vad det betyder .
Resolutionen begär parallellt nya medbeslutandebefogenheter för Europaparlamentet i fråga om invandring .
Man kan föreställa sig vad det kommer att göra av dem .
Såsom man kunde förutse har just Europeiska kommissionen gett parlamentet sitt stöd i det yttrande som den har avgett inför regeringskonferensen .
Vår grupp anser att det skulle vara mycket farligt att gå i den riktningen och att man tvärtom i dessa frågor måste stå nära folken och de nationella suveräniteterna .
Därför bör inte förfarandena i den första pelaren och förfarandena för den inre marknaden införlivas på identiskt sätt på områdena för säkerhet , rättvisa och utrikespolitik .
När det gäller dessa områden måste regeringskonferensen hitta nya samarbetsförfaranden , inriktade på rådets politiska roll och en inomparlamentarisk kontroll som utövas av de nationella parlamenten .
( Applåder ) Herr talman !
Jag talar som företrädare för den spanska delegationen av Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater , för delegationen av det spanska folkpartiet , beträffande Terrón i Cusís resolution om området med frihet , säkerhet och rättvisa .
Faktum är att vi inte i alla omröstningar har följt direktiven från Europeiska folkpartiets grupp , och vi har röstat för Terrón i Cusís resolution som på det hela taget är en utmärkt resolution .
Däremot röstade vi emot punkterna 2 och 6 , för vi anser att de är oriktiga juridiskt sett .
I stället har vi röstat för skäl J som ligger i linje som det jag själv , som föredragande av yttrandet , har föreslagit utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikesfrågor inför regeringskonferensen .
Vi har likaså röstat för punkt 13 .
En ändamålsenlig stadga och fri rörlighet och etablering för tredje land är något som det spanska folkpartiet länge har försvarat .
Av liknande skäl har vi röstat för punkt 14 där , i och med det muntliga ändringsförslaget en viss , högst berättigad oro för problem med subsidiariteten har beaktats , och där både vad gäller de politiska rättigheterna , inte längre rösterna i kommunvalen , utan de politiska rättigheterna i generella termer , ingår i medlemsstaternas suveränitet .
I och med det muntliga ändringsförslaget tyckte vi att vi kunde rösta för detta och det har vi också gjort . .
( DA ) De danska socialdemokratiska ledamöterna av Europaparlamentet har valt att rösta för resolutionsförslaget , men betonar samtidigt att vissa områden strider mot det undantag som Danmark har på det rättsliga området - ett undantag som den danska delegationen i PSE-gruppen naturligtvis vill respektera . .
( FR ) Detta betänkande , som jag inte har röstat för , handlar i mindre grad om mänskliga rättigheter än om " gemenskapsinförlivande " , i själva verket konsolideringen av fortet Europa .
De " framsteg " från 1999 som tas upp i betänkandet är bara framsteg i förhållande till Dublinkonventionerna och Schengenavtalen , och ännu en handlingsplan från Tammerfors , som inskränker invandrarnas rättigheter .
För i förhållande till mänskliga rättigheter är det en tillbakagång .
Europa fortsätter att avvisa personer till länder som anses farliga av FN : s flyktingkommissariat medan en del länder i Central- och Östeuropa som är EU-kandidater tar emot zigenarflyktingar som i mängd avvisats från Belgien .
Albaner från Kosovo och serbiska desertörer förvägras flyktingstatus medan Pinochet i lugn och ro klarar sig undan sin process .
Schengenkonventionens Europa jagar avgjort lättare förföljda från söder än diktatorer , samtidigt som FN anser att vi kommer att behöva 159 miljoner invandrare för att behålla den demografiska balansen från och med nu till år 2025 .
Europa bör legalisera alla personer som är utan uppehållstillstånd , ge dem asylrätt och rösträtt till alla val och sedan kan vi i kammaren tala om ett område för frihet och rättvisa .
Betänkande ( A5-0026 / 2000 ) av McCarthy Herr talman !
Jag vill börja med att påpeka att jag som borgmästare i Bilbao på nittiotalet fick tillfälle att lägga fram ett av de första urbana pilotprojekt som kommissionen skulle ge anslag till .
Våra erfarenheter i Bilbao av detta pilotprojekt har lett fram till fyra slutsatser : den första är att Europa måste behålla en urban politik och , i stället för att minska resurserna från 900 miljoner euro under föregående femårsperiod till 700 för innevarande femårsperiod , bör öka finansieringen av programmet , till exempel - så som vi i Gruppen De gröna / Europeiska fria alliansen har föreslagit - genom att i Urban-projekten åter investera den del av strukturfonderna som varje medlemsstat inte har förbrukat inom fastställt datum .
För det andra bör insatserna , när det är dags att besluta vilka områden man bör ge anslag till , koncentreras till projekt med en genomgripande verkan .
Spridda åtgärder är inte effektiva .
Man måste välja , och prioritera de värsta och mest överhängande fallen , till förmån för de fasta målen i sin helhet , det vill säga för de sociala , ekonomiska och miljömässiga aspekterna med en demokratisk förvaltning , liksom förhållandet mellan dem .
För det tredje bör man ta hänsyn till den synergism som ger upphov till andra gemenskapsprogram , liksom möjligheterna till en hållbar utveckling inom den miljö eller det område som avses .
Slutligen måste man lita på de instanser som finns närmast medborgarna , nämligen kommunerna och de lokala organen och stödja dessa .
Det är främst där man känner till de sociala behoven , där man är starkast engagerad i problemen och dessutom där man kan föreslå projekt och genomdriva dem på ett effektivt sätt utan att belasta dem med byråkrati och uppnå de bästa resultaten .
Slutligen , av våra fyra ändringsförslag i dagens omröstning har två antagits medan de övriga två förkastades .
Det tvingar oss att avstå i den slutgiltiga omröstningen , för vi inser inte varför inte miljöaspekten beaktas när det att dags att fatta beslut om vilka projekt som skall finansieras , och vi begriper inte varför man inte godtar att varje medlemsstat kan avsätta den del av strukturfonderna till Urban-projekten som de inte har förbrukat i enlighet med gemenskapsprogrammen .
Herr talman !
Jag skulle vilja påminna om att vi har haft många diskussioner i utskottet för regionalpolitik , transport och turism om Urban-initiativet .
Många idéer har framförts .
Jag skulle också vilja påminna om att det trots allt var det minsta gemenskapsinitiativet som fanns och att vi följaktligen hade föreslagit att anslaget skulle ökas genom ett ändringsförslag , som förkastades .
Vi beklagar detta eftersom det nämligen fanns kvar pengar från strukturfonderna i en del länder och dessa pengar skulle verkligen ha kunnat stödja pilotprojekt , eftersom Urban-projekten , vill jag påminna om , just är pilotprojekt som gör det möjligt att genomföra en verklig politik för städerna .
Jag skulle också här vilja uppmärksamma kommissionen på sammanhållningen mellan de olika politikområden som genomförts och jag skulle också vilja att kommissionen gör en sammanhållning av Urban-projekten med de framtida projekten från den budgetpost som kallas " hållbar stadspolitik " .
Herr talman !
Jag skulle slutligen också vilja påminna om att vi i dag fortfarande inte har någon europeisk politik för städerna i Europeiska unionen och jag vill klargöra att denna punkt , kanske , skulle kunna utvidgas inom ramen för omorganisationen och regeringskonferensen så att Europeiska unionen äntligen också får en verklig politik för städer .
Herr talman !
Jag skulle vilja påpeka att jag röstade för detta betänkande om hållbar stadsutveckling , vid namn Urban .
Liksom alla de andra gemenskapsinitiativen är det någonting mycket positivt .
Europa visar sig närvarande just i det ögonblick när man gör någonting för alla europeiska medborgare och inte bara för en enskild stads utveckling , vilken det vara må .
Med Urban vill man hitta lösningar på städernas förfall , och detta är någonting som intresserar de äldre mycket och som därmed intresserar Pensionärspartiet mycket .
Det finns ingen som har det sämre än en äldre människa i staden .
Jag hoppas att detta gemenskapsinitiativ kommer att bli ett föredöme för hur man löser problemet med äldre i städerna . .
( DA ) Vänsterns fem ledamöter av Europaparlamentet har valt att stödja Leader + , Equal-initiativet och Interreg , men inte Urban .
Vid en kommande granskning av dessa program bör EU : s insats koncentreras på gränsöverskridande uppgifter och anpassas till en utvidgning av EU .
Vi har röstat för betänkandet om meddelandet från kommissionen om fastställande av riktlinjer för ett gemenskapsinitiativ för ekonomisk och social förnyelse av städer och förorter som befinner sig på tillbakagång för att främja en hållbar stadsutveckling ( Urban ) .
I grunden är vi emot denna typ av program och strukturfonder , men eftersom omröstningen endast behandlar hur - och inte om - dessa resurser skall användas , har vi endast tagit ställning till innehållet och anser allmänt att förslaget om förnyelse av städer och förorter som befinner sig på tillbakagång innehåller förnuftiga slutsatser samt goda förslag och kriterier för projekten . .
( FR ) I betänkandet räknas allmänna begrepp upp rörande vad som kallas en strategi för urban förnyelse av stadskärnor och förorter som drabbats av den kapitalistiska ekonomins kris och dess konsekvenser : ökad arbetslöshet , utestängning och ungdomsbrottslighet .
I betänkandet understryks att för att säkra en hållbar utveckling i städerna , gäller det att genomföra en urban politik som inte åsidosätter de främsta offren för den ekonomiska krisen : arbetslösa , invandrare , flyktingar , kvinnor och utestängda .
Men det sägs ingenting om skälen och de ansvariga till krisen .
I betänkandet är det bara i bästa fall fråga om att rätta till vissa aspekter och efterverkningar av den .
Och dessutom med chockerande neddragna medel , eftersom enligt betänkandet själv är anslagen som tilldelats programmet Urban II för perioden 2000-2006 omkring 30 procent lägre än anslagen från den föregående perioden , som redan var låga ( 900 miljoner euro ) trots att det handlar om ett femtiotal projekt i hela Europa , vilket är obetydligt , när det är strängt taget samtliga storstadsförorter i vår världsdel och rentav stadskärnor som drabbas .
Därför röstar vi regelbundet för de konkreta åtgärder som anmälts för att hjälpa de minst gynnade sociala kategorierna , men vi avstår i fråga om själva betänkandet genom att ange att det härrör från fromma önskningar som finansierats med rabatt . .
( FR ) Fru föredragande , mina kära kolleger !
Jag måste säga att jag är mycket nöjd med att gemenskapsinitiativet Urban fortsätter , ett initiativ som siktar till att stödja den sociala och ekonomiska omvandlingen i städer och förorter i kris , detta för att främja en hållbar utveckling i städerna .
Med omkring 80 procent av den europeiska befolkningen boende i stadsmiljö är städerna i centrum av den ekonomiska , sociala och kulturella utvecklingen i Europa .
Samtidigt är de sociala och ekonomiska problem som det europeiska samhället brottas med mer markanta i städerna .
Många europeiska städer har nämligen en intern regional brytning : samexistensen , i städerna , av kvarter där man bedriver verksamheter med högt mervärde och där höginkomsttagare är bosatta och av kvarter , som markeras av låga inkomster , hög arbetslöshet , medelmåttiga och överbefolkade bostäder och ett starkt beroende av socialstöd .
Koncentrationen av sociala och ekonomiska problem till vissa stadsområden kräver en målinriktad intervention som tar hänsyn till problemens komplexitet .
Därför har Europaparlamentet krävt och lyckats uppnå en förlängning av gemenskapsinitiativet Urban i reformen av strukturfonderna .
Urbans framgång under programplaneringsperioden 1994-1999 är obestridlig .
Resultatet är påtagligt när det gäller förbättring av livskvaliteten i de målinriktade områdena .
Detta gemenskapsinitiativ främjade utvecklingen av goda metoder inom de ekonomiska , sociala och miljömässiga sektorerna .
Det hade dessutom fördelen att stärka rollen för de lokala myndigheternas , icke-regeringssektorns och de lokala myndigheternas roll och främja nya partnerskapsformer på området förförnyelse av städer .
Med det nya initiativet skall vi fortsätta att försöka nå dessa mål genom att stärka dem samtidigt som vi särskilt tar hänsyn till främjandet av lika möjligheter för män och kvinnor och integrationen av kategorier av människor som är socialt marginaliserade och missgynnade .
Vi kan således glädja oss åt att det antagits .
Man måste emellertid medge att på det finansiella planet kan vi inte utropa segern !
Det avsatta finansiella totalanslaget är nämligen inte på långa vägar i nivå med det som står på spel .
Anslagsbeloppet var 900 miljoner euro för perioden 1994-1999 och det är 700 miljoner euro för perioden 2000-2006 , det vill säga en minskning med 30 procent !
Denna minskning av finansmedlen har lett till en minskning av antalet program inom ramen för det nya Urban-initiativet .
Det valda taket tycks vara för lågt .
Det har satts till femtio projekt .
Det bör således ökas för att regionala och lokala faktorer skall beaktas samtidigt som de finansiella anslagen avsedda för medlemsstaterna behålls .
Mot bakgrund av denna koncentration på ett antal begränsade projekt spelar kanske offentliggörande och spridning av resultaten från det nya gemenskapsinitiativet Urban en viktig roll för att få en ökningseffekt .
På förslag av kommissionen minskades antalet städer som kan dra nytta av det nya Urban-initiativet för perioden 2000-2006 från 100 till 50 samtidigt som anslagen minskades med 30 procent .
Förslaget är till stort förfång för Portugal , trots att det är det land inom Europeiska unionen som har störst brister på det här området .
Man har gått ned till knappt två finansierade projekt , medan man för Tyskland räknar med tio , för Förenade kungariket nio och för Italien åtta .
Nåväl , fram tills nu har Portugal fått sex projekt finansierade , vilket har gynnat kommunerna i Porto , Gondomar , Lissabon , Odivelas , Oeiras och Amadora .
Det är därför absolut nödvändigt att kommissionen ser över sin ståndpunkt igen , särskilt beträffande tilldelningen av projekt till Portugal , så att förutsättningar skapas för att gå vidare och väcka liv i det ekonomiska och sociala arbetet i städer och förorter så att en hållbar tillväxt kan garanteras . .
( FR ) Betänkandet McCarthy om gemenskapsinitiativet Urban ger oss tillfälle att diskutera om det är lämpligt att gemenskapen ingriper på stadsområdet .
Situationen i vissa stadsområden är alarmerande och den sociala nöden visar sig i form av arbetslöshet , fattigdom och kriminalitet .
Narkotikahandeln i synnerhet underhåller osäkerhet och småbrottslighet .
Strukturfondernas effektivitet är tvivelaktig inför sådana sociala utmaningar .
Subsidiariteten borde leda till att vi erkänner att staten i utövandet av sina regeringsfunktioner och de lokala myndigheterna är mest lämpade för att ingripa på rätt sätt , staten genom att trygga den allmänna säkerheten och de lokala myndigheterna genom att hjälpa människor i svårigheter .
Även om man kan glädja sig åt viljan att skapa ett system för utbyte om lyckade företag , kan man inte ställa de specifika problemen för varje stadsområde på samma plan .
Gemenskapsinitiativet Urban ingår i Europeiska unionens vilja att införliva stadspolitiken i gemenskapen .
Det skulle vara mera relevant om Europeiska unionen inriktade sina finansiella ansträngningar på redan befintliga europeiska politikområden .
En del grupper och personer passar självklart på tillfället att ge sig in på ett nytt budgetöverbud , ett överbud som är speciellt illa valt vid en tidpunkt då staternas budget tvingas till en allvarlig avmagringskur på grund av EMU : s konvergenskriterier .
McCarthy föreslår således en ökning av de avsatta anslagen till Urban och främjande av detta gemenskapsinitiativ genom en dyrbar kommunikationskampanj som kommer att användas till att berömma det federala Europas goda gärningar .
Måste man påminna om att en utgifts effektivitet inte mäts i storleken på de anslag som tilldelas projektet ?
Däremot anser mottagarna av alltför många och höga subventioner att dessa på sikt kan tas för givna .
Målsättningen bör inte vara att stödja medborgarna utan att få dem att ta ansvar .
I betänkandet betonas slutligen starkt åtgärder till förmån för etniska och sociologiska minoritetsgrupper .
Vi kan bara förkasta en minoritetspolitik som ofrånkomligen är farlig för den sociala sammanhållningen .
Å ena sidan , uppmuntras genom denna politik till integration av invandrare där det skulle vara nödvändigt att främja deras assimilering med mottagarlandets kultur för att undvika att etniska getton uppstår som blir en explosionsrisk i staden .
Å andra sidan , laborerar den med principen om positiv diskriminering , en politiskt korrekt illusion och minst lika skadlig , såsom den amerikanska presidenten har visat .
På grund av dessa orsaker kunde den franska delegationen i UEN-gruppen inte godkänna betänkandet McCarthy .
Betänkande ( A5-0028 / 2000 ) av Decourrière Herr talman !
Programmet Interreg ligger oss särskilt varmt om hjärtat .
Jag gläder mig liksom många av mina kolleger åt att parlamentet har kunnat behålla detta Interreg-initiativ .
Eftersom jag själv bor i området Sarre-Lorraine-Luxemburg i södra Belgien vet jag att det är där Europa skapas , där vi lever med Europa dagligen och medborgarna faktiskt ser till att den europeiska uppbyggnaden lever fullt ut .
Dessa förslag bör verkligen beaktas och hållbar utveckling bör redan införlivas i dem .
Varför påpekar jag det ?
Helt enkelt för att de förslag som nu läggs fram fortfarande alltför ofta är miljöförstörande , på det sätt som de läggs fram .
Att godkänna nya vägar , till exempel , det är att godkänna nya skadliga faktorer i Europeiska unionen och det går helt emot den politik , som vi föreslår , i fråga om kamp mot gasutsläpp med växthuseffekt , till exempel .
Jag ber också att kommissionen inom ramen för de projekt som läggs fram skall vaka över att miljöpelaren i Europeiska unionens politik införlivas i dessa projekt och att målet att minska , till exempel , koldioxiden skall kunna vara ett pilotmervärde i de föreslagna projekten .
Jag tänker här särskilt på vissa infrastrukturer som håller på att genomföras .
Man vet att vissa medlemsstater fortfarande tvekar , till exempel , mellan järnväg och landsväg för genomfarter i känsliga områden såsom Pyrenéerna - jag tänker på Aspe-dalen .
Men jag tänker också på min region där min medlemsstat fortfarande tvekar mellan att bygga järnväg och en andra motorväg , A32 .
Sålunda också här ber jag således kommissionen att vara särskilt uppmärksam så att det blir en verklig sammanhållning mellan de olika politikområdena , i synnerhet i de framlagda Interreg-programmen .
Herr talman !
Jag röstade för Decourrières betänkande om gemenskapsinitiativet Interreg , framför allt på grund av det svar kommissionär Barnier gav några ledamöter som begärde att man i detta program skulle bry sig mer om de gränsregioner som har havsgränser .
Detta gjorde jag inte bara för att jag är född i en kuststad , Genua , utan framför allt för att även de gränser som utgörs av vatten är gränser .
Dessa gränser vetter mot Afrikas länder och Mellanöstern : vi måste ta större hänsyn till det faktum att det är viktigt att utveckla också kustregionerna i alla delar av Europa . .
( FR ) I min egenskap av ledamot av Europaparlamentet från ett gränsområde emotser jag med stort intresse det tredje Interreg-initiativet .
Vi kan aldrig tillräckligt påminna om de svårigheter som fanns förr i tiden i de områden vid gränserna , på land eller till havs , som hade delats ekonomiskt , socialt och kulturellt .
På grund av närvaron av gränser omvandlades de till yttersta randområden i de stater där de ingick , vilket alltför ofta ledde till att de statliga myndigheterna åsidosatte dessa områden inom ramen för den nationella politiken .
Därför infördes gemenskapsinitiativet Interreg från och med 1990 .
Syftet med programmet var att uppmuntra till gränsöverskridande , transnationellt och interregionalt samarbete samt en balanserad utveckling av gemenskapens område för att stärka den ekonomiska och sociala sammanhållningen i unionen .
Interreg syftar huvudsakligen till att finansiera gemensamma metoder för utveckling av små och medelstora företag , yrkesutbildning , grundutbildning , kulturellt utbyte , hälsofrågor , miljöskydd och miljöförbättring , kraftnät , transport och telekommunikationer .
Jag vill framhålla att det interregionala samarbetet bidrar till att ansluta de lokala och regionala myndigheterna till den europeiska integrationsprocessen .
Vi måste nämligen främja ett aktivare deltagande av de lokala och regionala myndigheterna när det gäller gemenskapsinitiativen , samtidigt som vi tar hänsyn till att de regionala och lokala myndigheterna ofta har mycket begränsad samarbetskapacitet på grund av mångfaldiga rättsliga ramar och utvecklingsnivåer på ena eller andra sidan av samma gräns .
Inom ramen för det gränsöverskridande samarbetet bör vi lägga större vikt vid att förbättra driftsvillkoren för sysselsättningsskapande små och medelstora företag .
På samma sätt och mot bakgrund av att femtio procent av arbetslösheten är strukturell arbetslöshet bör de medel som ställs till förfogande från Interreg vara tillräckligt stora för att komplettera nationella sysselsättningsfrämjande åtgärder .
Mer konkret kan sägas att den gränsöverskridande rörligheten omöjliggörs , bromsas och blir problematisk på grund av hinder , som alltför ofta är anknutna till skattesystemet ( dubbelbeskattning ) och det sociala trygghetssystemet .
Jag önskar att de projekt som ingår i programmen skall bidra till att finna lösningar på dessa problem och ge ett konkret innehåll åt den fria rörligheten för arbetstagare , en princip som i min region väger tungt !
Interreg-anslagen bör också bidra till att inrätta ett europeiskt forskningsområde .
Slutligen och framför allt finns det mycket stora förväntningar i regionerna på detta initiativ , eftersom kommunerna som inte är stödberättigade till mål 2 hoppas bli kompenserade tack vare Interreg !
Det är således viktiga saker som står på spel : införlivandet av gränsområdena kommer att utgöra en väsentlig faktor när den framtida europeiska regionalplaneringspolitiken utarbetas !
Jag hoppas att var och en är lika medveten om det som F. Decourrière som jag gratulerar ! .
( FR ) Gemenskapsinitiativet Interreg är en olycksdiger beståndsdel i den europeiska regionalpolitiken .
Denna politik som till ytan verkar generös eftersom den officiellt är avsedd för att hjälpa områden i svårigheter är en narrarnas marknad för de franska skattebetalarna .
Frankrike som bidrar med 17 procent av den europeiska budgeten , får bara 8 procent av de regionala strukturfonderna .
Mellan 1994 och 1999 fick våra regioner genomsnittligen 15,4 miljarder franc per år , men de kommer bara att få 14,7 miljarder mellan åren 2000 och 2006 .
Min region , Nord-Pas-de-Calais , kommer att särskilt beröras , eftersom franska Hainaut förlorar mål 1-stöden .
En oberättigad indragning i ett område vars främsta verksamheter har förstörts genom frihandelspolitiken i Europa .
Den europeiska regionalpolitiken stärker också Bryssels centralregering , med vilken de regionala myndigheterna uppmanas förhandla direkt om användningen av strukturfonderna .
Det är regionernas Europa , regioner som inte har samma kraft som våra nationer och lätt kommer att foga sig efter Bryssel .
Interreg-initiativet som tillkom 1990 för att förbereda - jag citerar : " gränsområdena till ett Europa utan gränser , således utan nationer , passar mycket väl in i denna filosofi " .
Decourrière framför emellertid kloka reflexioner då han pekar på Brysselteknokraternas brister .
Dessa kommer i synnerhet att leda till ett försenat genomförande av Interreg III och således finansiella förluster för mottagarområdena .
Vi är också ense med honom om att begära mer uppmärksamhet åt små och medelstora företag och naturligtvis vägra ta hjälp av ett externt tjänsteföretag .
Det är sådana metoder som ligger bakom den föregående kommissionens korruptionsaffärer .
Dessa punkter , som innehåller sunt förnuft och som vi har röstat för , rättar dock inte till den eurofederalistiska filosofi som präglar gemenskapsinitiativen , i synnerhet Interreg .
Därför röstade Nationella fronten emot betänkandet . .
( FR ) Europaparlamentet har gett sin åsikt om kommissionens riktlinjer rörande gemenskapsinitiativet Interreg om gränsöverskridande , transnationellt och interregionalt samarbete .
Jag vill försvara ett ändringsförslag som ingavs av min grupp om frågan om detta initiativs havsdimension .
Det handlar inte om att åter oroa sig för Atlantbågens framtid utan om nödvändigheten att införliva principen om havsgränser i avdelning A rörande det gränsöverskridande samarbetet .
I Europeiska kommissionens riktlinjer finns det inte många havsområden som är stödberättigade till Interreg III A. Ändringsförslagen till betänkandet Decourrière går mot en " havsinriktning " av Interreg .
Denna utveckling är viktig och bör fortsätta eftersom det är unionens framtid som står på spel .
Jag känner till Europeiska kommissionens motstånd i frågan .
Den framförde det vid samtalet i november om framläggandet av Interreg III .
Men jag vill påpeka följande : att förhindra ett erkännande av havsgränserna betyder att man förnekar att det finns ett område som är potentiellt rikt på projekt och innovationer .
Ett enda exempel : det så kallade " keltiska " området som omfattar områdena Bretagne i Frankrike , Cornwall och Devon i Förenade kungariket , Cork och Waterfold i Irland är ett område som har en närekonomi grundad på beroende av fiskerisektorn och betydelsen av lantbruket samt privilegierade kulturella och vänskapliga band ( vänorter ) .
Interreg III , avdelning A , skulle göra det möjligt för dessa områden att föra fram ett antal strukturprojekt som är nödvändiga för utvecklingen av små och medelstora företag samt för teknisk forskning och utveckling genom kunskapsöverföring .
Det skulle således vara önskvärt att Europeiska kommissionen kan delta i genomförandet av infrastrukturer för hamnar och flygplatser för förbindelserna mellan regionerna .
Denna politik skulle således få stora ekonomiska konsekvenser för fisket i Bretagne eftersom fisken skulle kunna landsättas på framskjutna irländska baser för att därefter skickas hem till livsmedelsföretagen i Bretagne .
Införandet av havsgränsen i avdelning A skulle göra det möjligt att äntligen erkänna ett enda ekonomiskt och stort område i västra randområdet inför Europeiska unionens kontinentala förskjutning .
Det skulle vara att visa respekt för dessa yttersta randområden som oroar sig en aning inför utvidgningen mot öster .
Havsvärlden har en stor potential .
Vi får inte åsidosätta den i gemenskapens nydanande pilotprogram som gör det möjligt att fastställa Europas nya geografiska och ekonomiska karta . .
( DA ) Det europeiska projektet startade som ett samarbete mellan stater .
Detta samarbete har säkrat freden och stabiliteten i vår del av Europa i över 50 år .
Som ett resultat av de ekonomiska och politiska framgångarna i vår del av världen , som bl.a.
EU är ett bevis på , och i och med den allt större spridningen av våra västliga värderingar , har konkurrensen på världsmarknaden vuxit kraftigt under de senaste årtiondena .
Denna konkurrens skall EU vara redo att möta .
Det kan vi bara göra genom att intensifiera samarbetet inom gemenskapen .
Här handlar det inte om en större integration av länderna i form av en federation , utan om att utnyttja våra ekonomiska möjligheter över gränserna .
Projekt som gör det möjligt att bygga ekonomiska tillväxtcentrum på gemenskapsnivå , som kommer att kunna anta utmaningen från våra konkurrenter på det globala planet .
Jag välkomnar därför en fortsättning på programmet . .
( FR ) Betänkandet av Decourrière saknar inte goda egenskaper ; denna lika tydliga som uttömmande presentation av Interreg-initiativet och dess roll för att bryta gränsregionernas isolering ställer sig , i punkt 16 , på de små och medelstora företagens sida .
Med min kollega Dominique Souchet , som är insatt i denna fråga , har jag ingivit fem ändringsförslag som framhåller de små och medelstora företagens och hantverkarnas roll inom ramen för Interreg , betydelsen av samarbete mellan företag och kravet på att ekonomiska och sociala partner skall vara delaktiga i utformningen och genomförandet av programmen .
Dessa ändringsförslag har antagits enhälligt , vilket gläder mig .
Men den franska delegationen i vår grupp kan inte acceptera att kommissionen och den federalistiska klanen avleder Interreg-initiativet från dess syfte , för att ytterligare försvaga nationernas politiska roll .
Vi avser inte att låta Bryssel ta hand om medlemsstaternas regionala fysiska planering , vilket skäl L i betänkandet antyder .
Vi begär bara en sak från kommissionen : att den nöjer sig med att se till att genomförandet av gemenskapens politik inte hotar en balanserad fysisk planering .
Den gemensamma jordbrukspolitiken och EMU : s skadliga effekter för balansen mellan olika regioner och framför allt för vitaliteten i de mest avlägsna och glesbefolkade landsbygdsregionerna , visar att en sådan ambition är allt annat än ett latmansgöra .
Därför kan vi inte godkänna utvecklingen av området IIIC i gemenskapens initiativ , ett område som genom att uppmuntra samarbetet mellan regionerna under kommissionens ansvar håller medlemsstaterna vid sidan om .
Den förtjusning som uttrycks för område IIIC blir desto märkligare då föredraganden i sin motivering själv erkänner att " utkastet till riktlinjer [ innehåller ] inga uppgifter om eventuella samarbetsområden " ( s.16 ) och att " ansvaret är [ ... ] oklart " ( p.17 ) .
Att under sådana omständigheter kräva ytterligare medel för detta avsnitt , som i punkt 20 , är ännu ett av de lika oansvariga som ideologiska överbud som kammaren är sin vana trogen .
Låt oss till sist konstatera det felaktiga i den vilja som uttrycks såväl i kommissionens dokument som i betänkandet av Decourrière : att Interreg skulle användas för freden och återuppbyggnaden på Balkan .
Jag tror inte att strukturfonderna skall utnyttjas för att reparera de skador som amerikanerna har åsamkat Serbien i samband med de både brottsliga och ineffektiva bombningarna .
Det är Washingtons sak och inte vår , att ta på sig ansvaret för en konflikt som de utlöste för att tjäna sina egna intressen .
Därför har den franska delegationen i vår grupp inte kunnat stödja Decourrièrebetänkandet .
Vi har valt att avstå vid den slutliga omröstningen .
Betänkande ( A5-0025 / 2000 ) av Procacci Herr talman !
Jag röstade för Procaccis betänkande om landsbygdsutveckling , inte bara för att jag instämmer i huvuddragen i Leader-programmet utan också för att det är den andra sidan av Urban-programmet , som vi talade om tidigare .
Precis som de äldre i städerna är mycket ensamma börjar de äldre på landsbygden bli den enda kvarvarande befolkningen , eftersom de unga flyttar till städerna : de dras till ljusen , till barerna också , och landsbygden töms .
Jag tror alltså att det är mycket viktigt att detta projekt inom Europeiska unionen får stöd av alla och byggs ut ytterligare .
Herr talman !
Jag är angelägen om att här hänvisa till en aspekt , som i stor utsträckning försummades i gårdagens debatt när det gäller programmet Leader + , som förhoppningsvis snart skall påbörjas .
Men framför allt vill jag också utnyttja tillfället att uttrycka mitt fullständiga godkännande av tyngdpunkterna i kommissionens nya program .
Detta gäller i synnerhet för det integrerade förfarandet med flera sektorer , vilket ökar allt mer i betydelse när det gäller jordbruket och som också alltid framhävs av jordbruksministrarna i medlemsstaterna .
Men även det faktum att man lägger mer vikt vid miljöskyddet när det gäller landsbygdsfrågor är av stor betydelse för allas vår framtid .
Att jordbrukarna kallas för förvaltare av landsbygden ger väl bäst uttryck för vilken riktning den kommande jordbrukspolitiken i ökande utsträckning tar , och naturligtvis genomförandet av den .
Jag anser också att det är mycket positivt att en av de väsentliga ändringarna av Leader + -programmet består i att nu all landsbygd och därigenom 80 procent av EU : s totala yta , respektive 25 procent av befolkningen i de 15 medlemsstaterna , kan dra nytta av programmet .
Ändå har det totala anslaget om 2 020 miljoner euro för sexårsperioden satts lågt , ja alltför lågt .
Dessutom , och det är framför allt det jag också anser att det handlar om , har man ännu inte räknat med några specifika initiativ för bergsområdena .
Inom ramen för Leader + -programmet refererar parlamentet till glesbygdsområdena i Nordeuropa , men inte till de lika ofta mycket glest bebyggda och därigenom missgynnade bergsområdena .
Tack för er uppmärksamhet ! .
( PT ) Det gemensamma initiativet Leader + , även om det är en fortsättning på tidigare initiativ , uppvisar en del besynnerligheter .
Först och främst halveringen av de tillgängliga anslagen , trots att perioden förlängts .
Likväl inkluderas nya mål , till exempel finansieringen av Natura nätverk 2000 , och landsbygden blir ett annat valbart alternativ .
Trots att det här gemenskapsinitiativet avser landsbygdens tillväxt tar man inte samstämmigt upp jordbruket och jordbruksproduktionen , och detta är inte rimligt .
Ingen landsbygd utan jordbruk , vilket gör att vilken strategi som helst för landsbygdens tillväxt måste baseras på jordbrukets endogena potential , oaktat andra aktiviteters större eller mindre tillväxt för att hindra landsbygdens desertering .
Därför menade vi att det var så viktigt att förbättra betänkandet med de förslag som vi lade fram om att jordbruksaktiviteterna och lantbrukarna uttryckligen borde inkluderas i strategin för landsbygdens tillväxt , och att man borde ansöka om större anslag så att man kan fortsätt med programmet på de orter som tidigare inkluderats samt ta det nya programmet , som skall fortsätta att privilegiera de minst gynnade områdena , i försvar .
Min inställning till Leader hänger samman med min inställning till EU : s jordbrukspolitik över huvud taget .
Såväl Leader I som Leader II , vilka genomförts under 1990-talet , har ingått i den nya gemensamma jordbrukspolitik som tillämpats allt sedan revideringen 1992 och har tillsammans med andra åtgärder utgjort den s.k. andra pelaren i EU : s politik för landsbygdsutveckling .
Deras verkliga syfte har varit att förringa och skyla över de katastrofala följderna av den nya gemensamma jordbrukspolitiken och att vilseleda de små och medelstora jordbruken , och de har inte haft till syfte att utveckla landsbygden och att behålla jordbruksbefolkningen på landsbygden , vilket man så hycklande brukar påstå .
Detta framgår av det faktum att jordbruksinkomsterna och sysselsättningen har minskat mycket hastigt i de områden där dessa initiativ har tillämpats , vilket lett till allt snabbare avfolkning av dessa områden .
Grekland är ett betecknande exempel .
Som mål 1-land omfattades Grekland i sin helhet av gemenskapsinitiativen från Leader .
Samtidigt minskade sysselsättningen inom jordbruket med 2,3 procent under perioden 1994-1999 , medan jordbruksinkomsterna minskade med 15,2 procent .
Jag anser att Leader + kommer att vara effektivare än Leader I och II av följande orsaker .
De verkliga målen för Leader + är de samma som för Leader I och II .
Dvs. att mildra och skyla över de negativa effekterna av den gemensamma jordbrukspolitik som kommer att tillämpas inom ramen för Agenda 2000 .
Men denna gemensamma jordbrukspolitik är sämre än den föregående och dessutom har den ett sämre utgångsläge , eftersom revisionen av den gemensamma jordbrukspolitiken 1992 och GATT-avtalet 1995 har lett till betydande problem och svårigheter för jordbruksekonomin .
Urvalskriterierna och de verksamheter som finansieras genom Leader kan i bästa fall lindra enstaka mindre viktiga landsbygdsproblem , men i värsta fall urartar de till offentliga utgifter som bara tjänar till att döva samvetet .
Programmen leder inte till någon allsidig utveckling av de utvalda områdena och de leder inte heller till nya , stadigvarande arbeten på landsbygden , för de flesta verksamheterna har inte någon produktiv inriktning .
De verkliga anslagen till Leader + är mindre än anslagen till Leader II , trots en ökning med 15 procent ( från 1775 miljoner euro för Leader II till 2020 miljoner euro för Leader + ) .
Och detta beror på att ökningen med 15 procent är nominell och inte reell , eftersom den genomsnittliga årliga inflationen inom gemenskapen under dessa år uppgår till ungefär 2 procent .
Leader + pågår ett år längre än Leader II .
Till Leader + kan man föra alla EU : s regioner , medan Leader II omfattade mål 1-regionerna och vissa regioner inom mål 5b och 6 .
Men jag vill påpeka att även om de reella anslagen till Leader + var högre , så skulle gemenskapsinitiativet ändå vara ineffektivt , eftersom den jordbrukarfientliga inriktningen av den gemensamma jordbrukspolitiken inom ramen för " Agenda 2000 " inte kan vare sig kompenseras eller mildras av sådana program som i många områden endast syftar till att skyla över , att vilseleda och att döva samvetet .
Jag motsätter mig många av åsikterna i betänkandet .
Jag vill ännu en gång påpeka de negativa förändringarna i den gemensamma jordbrukspolitiken ( 1992 - Agenda 2000 ) .
Jag anser att Leader + inte kommer att bidra till en verklig lösning av landsbygdens problem , med allt svårare förhållanden för jordbruket , som ju har varit och bör vara den viktigaste samhällsekonomiska näringsgrenen på landsbygden .
Jag kommer för min del att informera jordbrukarna om syftet med dessa program .
Jag kommer att verka för att de skall utnyttjas på bästa tänkbara sätt utan att slösas bort och , framför allt , kommer jag att verka för att utveckla jordbrukarnas kamp mot den katastrofala gemensamma jordbrukspolitiken , som utarmar dem och leder dem till ekonomisk bankrutt , samtidigt som landsbygden avfolkas .
Om man inte avskaffar denna gemensamma jordbrukspolitik , finns det nämligen inget program som kan garantera att de små och medelstora jordbruken överlever och att landsbygden vitaliseras socialt och ekonomiskt . .
( FR ) Samtliga ledamöter i gruppen Unionen för nationernas Europa har röstat för nästan allt i betänkandet av vår kollega Procacci rörande gemenskapsinitiativet Leader + .
Vi har emellertid ändrat det förslag till betänkande som hade godkänts av utskottet för jordbruk för att klarlägga vissa punkter varvid gemenskapsinitiativet kunde göras mer operativt .
Det verkar för oss väsentligt att i synnerhet förenkla de administrativa och finansiella förfaranden som visade sig bli för tunga och långsamma inom ramen för initiativet Leader II .
Det verkar också nödvändigt att säkra att bättre hänsyn tas till de lokala aktörernas utvecklingsprioriteringar och att inte utdelningen av fonderna Leader + bara begränsas till jordbruksområden med låg befolkningstäthet .
I ändringsförslag 10 , som jag har ingett på min grupps vägnar , hänvisas till begreppet " ekonomisk och social sammanhållning " i stället för " regionalplanering " eftersom Europeiska unionen inte har erkänd befogenhet på området .
I ändringsförslag 11 ersätts termerna " statlig eller kommunal administration " med " samtliga offentliga förvaltningar " .
De lokala åtgärdsgrupperna bör visserligen utgöra en balanserad enhet som är representativ för partner från olika socioekonomiska miljöer i området men på beslutandeplanet bör i själva verket samtliga offentliga förvaltningar ( kommuner , län , regioner och stater ) företrädas i sin helhet vilket nivå de än har .
Föredragandens formulering var således alltför inskränkande , enligt vår åsikt .
Vad beträffar ändringsförslag 12 uppfyller det förväntningarna i Europaparlamentets utskott för regionalpolitik .
Det inbegriper den nödvändiga samordningen mellan Leader + och gemenskapsprogrammen för samarbete och partnerskap , såsom Interreg , Phare , Sapard eller Meda .
På Europeiska unionens , kandidatländernas och EFTA : s medlemsstaters territorium kan det finnas interna förbindelser mellan de olika gemenskapsinitiativen .
Man måste komma ihåg att de verkliga prioriteringarna för den europeiska världsdelen är att införa en operativ nivå inom europeisk ram och inte inom en global ram , såsom föredraganden föreslår .
Skapandet av organisationer liknande lokal åtgärdsgrupper ( GAL ) kan med fördel uppmuntras av Europeiska unionen , naturligtvis förutsatt att motsvarande kostnader bestrids av de olika parterna .
Vi ställer oss i grund och botten naturligtvis positiva till gemenskapsinitiativet Leader + .
Vi måste komma ihåg att vid konferensen om landsbygdsutveckling som hölls i Cork den 7-9 november 1996 definierades landsbygdsutveckling såsom en av Europeiska unionens prioriteringar eftersom det är av största vikt att bevara vårt jordbruks och hela landsbygdsstrukturens ( infrastrukturer , offentliga och privata tjänster ... ) integritet .
I det sammanhanget har vi i utskottet beklagat avsaknaden av anslag för landsbygdsutveckling och stött de ändringsförslag som begär en ökning av budgeten för detta gemenskapsinitiativ , så att det kommer i jämvikt med de tidigare initiativen Leader I och Leader II .
Jämfört med det senare initiativet som hade begränsad giltighetstid på sex år , är den anslagna budgeten för Leader + femtio procent lägre för en period av sju år .
Det är inte godtagbart med tanke på den betydande landsbygdsutvecklingen och konsekvenserna för jordbrukarna av pris- och stödsänkningarna enligt den planerade reformen av den gemensamma jordbrukspolitiken till följd av Berlinavtalen .
Bland de prioriterade kriterier som kommer att införas på europeisk nivå för att möjliggöra lokala anmälningar bör slutligen särskild uppmärksamhet ägnas åt de projekts kvalitet och originalitet som redan uppburits av GAL inom ramen för initiativet Leader II men som inte kunnat slutföras på grund av tidplanen och de omständliga planerade förvaltningsåtgärderna .
( Sammanträdet avbröts kl .
13.40 och återupptogs kl .
15.00 . )
 
Fodertillsatser Nästa punkt på föredragningslistan är betänkande ( A5-0015 / 2000 ) av Graefe zu Baringdorf för utskottet för jordbruk och landsbygdsutveckling om förslaget till rådets direktiv om ändring av direktiv 70 / 524 / EEG om fodertillsatser ( KOM ( 1999 ) 388 - C5-0134 / 1999 - 1999 / 0168 ( CNS ) ) . .
( DE ) Herr talman , kommissionär Byrne !
Direktiv 70 / 524 innebär nu en annorlunda behandling av de tekniskt högt utvecklade tillsatserna med tanke på ersättning av gällande tillstånd .
Här har nu kommissionen föreslagit att man skall genomföra en harmonisering i tillståndsförfarandet , så att de ämnen som godkänts före 1988 skall jämställas med dem som godkänns nu .
Så långt anser vi i utskottet för jordbruk och landsbygdens utveckling att allt är i sin ordning .
Men detta direktiv omfattar också godkännande av antibiotika , läkemedel , tillväxtbefrämjande medel och genetiskt modifierade organismer ( GMO ) .
Här handlar det om hälsa och inte om en enkel tillnärmning av rätten .
Därför anser vi i utskottet för jordbruk att den rättsliga grunden - artikel 37 - här inte kan godkännas , utan att kommissionen måste föreslå oss en rättslig grund i enlighet med artikel 152 , dvs. medbeslutande från parlamentet .
Vi har frågat utskottet för rättsliga frågor och den inre marknaden , som med tanke på denna tillnärmning av rätten har påpekat att artikel 37 skulle vara tillräcklig i detta fall .
Vi från utskottet för jordbruk har dock inte begränsat oss till behandlingen av denna tillnärmning av rätten , utan med tanke på att det i detta förslag också handlar om genetiskt modifierade organismer har vi lämnat in ytterligare ett ändringsförslag , och det går in på frågan om innehållet och därmed också på befolkningens hälsa .
Vi har i utsädesdirektivet förhandlat två år med kommissionen och kommit fram till en kompromiss , som i detta direktiv reglerar utsättningen av genetiskt modifierade organismer .
Vi har där utgått från den text som ligger till grund för detta direktiv 70 / 524 .
Vi kan inte förstå , herr Byrne , varför kommissionen , när den gör tillnärmningar , inte också gör en tillnärmning i texten som rör de genetiskt modifierade organismerna .
Vi har nu lämnat in ett ändringsförslag , som just behandlar ordalydelsen av denna kompromiss från kommissionen .
För övrigt har denna ordalydelse också övertagits i skogsodlingsdirektivet om användning av skogsodlingsmaterial , och vi anser att det är absolut nödvändigt att ta upp denna text nu också i detta direktiv .
Kommissionen har i utskottet hänvisat till att den har för avsikt att i framtiden lägga fram ett novel food-direktiv .
Detta bör dock inte vara något hinder för att man redan i detta fall företar en tillnärmning , så att det här inte uppstår någon rättslig osäkerhet beträffande olika direktiv .
Därför utgår vi från att ni också kommer att anta vårt ändringsförslag rörande dessa genetiskt modifierade organismer .
Det faktum att det fortfarande är den gamla texten som står i detta direktiv 70 / 524 har att göra med att utsädesdirektivet lades fram 1986 i parlamentet och att vi fram till 1988 förhandlade med kommissionen , medan betänkandet om detta direktiv behandlades 1994 , och uppenbarligen tillmätte då parlamentet inte de genetiskt modifierade organismerna samma betydelse som vi gjorde senare , när jag var föredragande .
Därför anser vi , kommissionär Byrne , att de ändringsförslag vi lämnat in bör antas av er även med avseende på den rättsliga grunden .
Om så inte är fallet , måste vi förbehålla oss rätten att återförvisa detta betänkande till utskottet , för att sedan , på liknande sätt som vi gjort beträffande utsädesdirektivet , förhandla med er om denna känsliga punkt , och här vill jag än en gång påpeka att den text som vi nu har utarbetat gäller som kompromiss både för er och för vår rättstjänst .
Vi måste alltså inte på nytt förhandla om texten , utan vi måste bara ta upp denna text i direktivet .
Jag är spänd på att få höra , kommissionär Byrne , vad ni kommer att säga om våra förslag !
( Applåder ) Herr talman , herr kommissionär !
Har regleringen av fodertillsatser att göra med konkurrens eller med konsumentpolitik ?
För kommissionen och utskottet för rättsliga frågor är det en fråga om konkurrens .
Säkerligen måste vi ta hänsyn till djurfoderindustrins konkurrenskraft när föreskrifterna för ämnen som tillåtits före och efter 1988 harmoniseras .
Det bör förhindras att priset på djurfoder höjs , och därför bör Doyles ändringsförslag 4 och 5 stödjas .
Men i första hand är det , som Graefe zu Baringdorf formulerat det i sitt betänkande , en konsumentpolitisk fråga .
Livsmedelssäkerheten måste ha absolut prioritet i alla diskussioner om djurfoder .
När vi talar om öppenheten i näringskedjan , så gäller det från dynggrepen till bordsgaffeln , och därför börjar alltså konsumentskyddet med djurfodret .
Antibiotika , tillväxtbefrämjande medel och genetiskt modifierade organismer hamnar ändå till slut i människans näringskedja .
Som en konsekvens av dioxinskandalen blev det klart för oss alla att vi äntligen måste ta oss ur detta mörka hörn .
Regleringen av fodertillsatserna är ett steg i rätt riktning .
Enligt artikel 152 i EG-fördraget är vi ålagda att undanröja sådana orsaker som kan hota människans hälsa .
Betoningen ligger entydigt på orsaker .
Helt konsekvent måste vi stänga av de ursprungliga källorna till skadliga ämnen - nämligen skadliga fodertillsatser .
I annat fall , anser jag , laborerar vi med symptomen , men vi bekämpar inte orsakerna .
Befolkningen är mycket kritisk i synnerhet när det gäller användning av GMO .
Vi måste ta hänsyn till befolkningens ökande känslighet beträffande GMO , och reglera användningen i djurfoder i enlighet med detta .
För det första : Om en tillsats består av genetiskt modifierade organismer , eller om den innehåller sådana organismer , får denna tillsats bara tillåtas om den är ofarlig för människans hälsa och för miljön .
För det andra : Det är förnuftigt att analogt med bestämmelserna i lagen om avyttring av utsäde , vilket även föredraganden har berört , utfärda föreskrifter för genetiskt modifierade fodertillsatser .
Och för det tredje : För att få en öppen konsumentpolitik behöver vi en märkning av genetiskt modifierat djurfoder .
Denna entydiga innehållsdeklaration för djurfoder möjliggör alltså en dubbel beslutandefrihet , både för den som använder djurfoder och för den senare konsumenten .
Beslutet bör ligga hos den myndigförklarade medborgaren , anser jag .
Vi talar alla om de skandalöst pungslagna medborgarna , som har förlorat förtroendet för livsmedelssäkerheten .
Med en konsekvent reglering av fodertillsatserna kan vi nu bidra väsentligt till att återvinna förtroendet .
Därför är jag alltså mycket spänd på att få höra ert svaromål vad gäller våra ändringsförslag .
Alltså kommer vi naturligtvis att rösta så att vi eventuellt skickar tillbaka förslaget till utskottet .
Herr talman , kära kolleger !
Föreliggande förslag till ändring av direktivet om fodertillsatser från år 1970 är det första i en hel rad förslag när det gäller djurfoder .
Vi kommer alltså under de närmaste månaderna här i parlamentet att diskutera ytterligare några .
Att denna fråga har central betydelse bevisar den stora uppmärksamhet som den europeiska allmänheten har skänkt skandalerna med dioxin , antibiotika , slam från reningsverk osv .
Det handlar här alltså om en viktig beståndsdel i skyddet av allmänhetens hälsa .
Därför anser vi att artikel 152 skall användas som rättslig grund och inte artikel 37 , som kommissionen har föreslagit .
Den ändring som kommissionen har föreslagit , nämligen lika behandling av de tillsatser som godkänts efter respektive före den 31 december 1987 , är oomtvistad , och har vårt fulla stöd .
Utskottet för jordbruk och landsbygdens utveckling har dock enhälligt gjort några viktiga ändringar i kommissionens förslag .
De av kommissionen föreslagna bestämmelserna medför risk för monopolbildning vid saluförandet av vissa tillsatser .
Förslagsrätt medges endast dem som erhållit det ursprungliga godkännandet , men utesluter de företag som senare har fått ett godkännande .
En sådan monopolbildning , som exempelvis skulle kunna leda till en höjning av priset på djurfoder , bör vi förhindra genom att ge ett preliminärt godkännande till alla företag som den 1 april 1998 saluförde ett visst ämne .
Detta skall sedan gälla tills den förnyade utvärderingen har avslutats .
Den viktigaste ändringen gentemot kommissionens förslag gäller dock det av föredraganden rekommenderade inkluderandet av bestämmelser om genetiskt modifierade organismer i direktivet om tillsatserna .
Han har här utgått från den kompromiss som parlamentet och kommissionen kommit överens om beträffande godkännande av genetiskt modifierade organismer utanför utsättningsdirektivet .
Denna utgör redan grundvalen för godkännandet av genetiskt modifierade organismer .
Därför är det bara logiskt och i enlighet med de bestämmelser som vi redan har godkänt på andra områden - jag kan bara nämna skogsodlingsmaterial - att även i föreliggande fall föreskriva bestämmelser om genetiskt modifierade fodertillsatser .
Här spelar i synnerhet märkningen av genetiskt modifierade tillsatser en viktig roll .
Å ena sidan medger den att jordbrukaren kan fatta ett medvetet beslut om huruvida han vill använda sådant djurfoder eller inte , och å andra sidan blir det möjligt för konsumenten att avvisa livsmedel som framställts på basis av genetiskt modifierade organismer .
Avslutningsvis också ett hjärtligt tack från vår grupp till föredraganden , som lagt ner mycket arbete på detta .
Jag tror vi kan vara nyfikna på att få höra vad Byrne kommer att säga .
Herr talman , ärade kolleger !
Detta betänkande handlar mer om formerna , dvs. hur tillsatsämnen skall godkännas , och något mindre om vilka de är och hur de fungerar .
Jag måste få ta tillfället i akt att understryka hur viktigt det är att alla dessa direktiv i fortsättningen behandlas enligt förfarandet i artikel 152 , eftersom både livsmedelssäkerhet och miljöfrågor kräver en sammanhållen politik , en helhetssyn .
Vi kan inte göra som vi gjort hittills , dvs. ta varje detalj för sig och ofta först när skadan redan är skedd .
Föredraganden har betonat prövning och märkning av GMO i fodertillsatsen .
Jag skulle än en gång vilja tala om antibiotika .
Förvisso är fem av de nio antibiotika som ursprungligen var tillåtna i foder i dag förbjudna , men det är oerhört viktigt att vi förbjuder även de sista fyra , inte bara för folkhälsans , utan även för djurens skull .
Vi har kommit så långt att vi känner till antibiotikaresistensens oerhörda hot mot folkhälsan , framför allt för småbarn .
I många medlemsstater kan man redan bevisa att missbruket i djurhållningen är helt onödigt .
Det finns flera länder som för länge sedan har fasat ut foderantibiotika , och det finns några som är på väg att göra det med lyckat resultat .
Försiktighetsprincipen , som vi talar mycket om , har vi för länge sedan gått förbi , när det handlar om antibiotika .
Det finns emellertid ytterligare en princip i miljöarbetet som är viktig , nämligen utbytesprincipen .
Jag skulle vilja säga något kort om coccidiostatika .
Det är ett tekniskt antibiotikum , som inte är absolut nödvändigt .
Det finns ersättningsmedel .
Det går att vaccinera kycklingar .
Det kostar visserligen litet mer , men är ofarligt för miljön .
I dag åker coccidiostatika ut med gödseln på åkern .
Därmed hamnar det i vattnet som ju faktiskt är vårt viktigaste livsmedel .
Herr talman , herr kommissionär , mina kära kolleger !
Betänkandet om fodertillsatser avser ett teknisk-ekonomiskt problem för att återställa konkurrensjämvikt mellan de olika fodertillsatserna och mellan tillsatsernas producenter .
Men nu efter den allvarliga dioxinkrisen som drabbade Belgien och andra europeiska länder förra sommaren kan man inte nöja sig med att diskutera om en enkel konkurrensfråga .
En gång i tiden , även om det gick mer obemärkt förbi allmänheten , upptäckte nämligen kommissionens vetenskapliga experter industriella kalkrester fulla med dioxin i pressade citrusfrukter som importerats från Brasilien .
Därför är det tid att redovisa samtliga beståndsdelar i den kedja som deltar i tillverkningen av foder för avkastningsdjur .
Vi kan i förbigående konstatera , och det är en skandal , att problemet är mycket mindre allvarligt när det gäller foder för våra hundar , katter och övriga husdjur .
Är det på grund av den vilda och globaliserade konkurrens som denna sektors industrier ägnar sig åt som den har omvandlats till en återvinningssektor för avfall från livsmedelssektorn ?
Ett så allvarligt ämne kan inte begränsas till en teknisk debatt även om det ju är det direktiv som begränsar tillståndet för antibiotika och andra tillväxtfaktorer .
De försiktighetsåtgärder som vi gör oss beredda att vidta för djurfoder bör också tillämpas i fråga om foder till lantdjur , just de djur som vi återfinner på tallriken .
Såsom det med kraft betonas i betänkandet är märkning en absolut nödvändighet så att varje jordbrukare i sitt företag känner till samtliga ingredienser som ingår i det foder som han avser att ge till sin besättning .
Han bör också veta om genetiskt modifierade organismer , GMO , har trängt in i hans proteinkornspåse .
Dessa beståndsdelar kan potentiellt utgöra en folkhälsorisk .
Genom försiktighetsprincipen har vi i varje fall fått krav om en tydligt angiven spårbarhet på alla nivåer vid saluföringen av dessa produkter .
Men före märkningen måste tydliga regler införas .
Man måste ställa enkla frågor såsom frågan om det verkliga syftet med användning av djurfoder .
Om vi betraktar alla problem som det har åsamkat oss ur etisk synpunkt och sanitär synpunkt , måste vi nu ställa oss frågan om själva användningen .
Det kapitel i vitboken om livsmedelssäkerhet , som behandlar djurfoder , bör i det avseendet tjäna som grund för arbetet med att gå långt bortom de enkla saluföringsfrågorna .
Kommissionen har vid flera tillfällen använt följande exempel : " från grepen till gaffeln " .
Vår kollega i PPE betonade det nyss .
Det är en god formulering , men vi måste också ge den mening .
Och för att ge den mening måste vi behandla såväl problemen med djuren som problemen med konsumenternas hälsa .
Därför är det viktigt att godkänna ändringsförslag 2 till skäl 4 , som gör det möjligt att undvika risk för monopol , om de bolag som först fick tillstånd att saluföra en tillsats skulle förbli de enda som kunde utnyttja det under omvärderingsperioden .
Men ändringsförslag 4 och 5 till den nya artikel 2 a måste framför allt godkännas , eftersom de gör det möjligt att tydligt utpeka tillsatser som är genetiskt modifierade för att användarna skall kunna fatta beslut med full sakkännedom .
Herr talman , mina damer och herrar ledamöter !
Användningen av tekniskt avancerade tillsatser inom djurfoderbranschen kräver detaljerad information från aktörerna - och det är som bekant ganska många - om deras insatser , för att man skall förhindra metoder som bryter mot gemenskapsrätten .
Det befintliga direktivet om fodertillsatser kan inte ensamt åstadkomma detta .
Det kommer att följas av andra direktiv , och jag anser att de är på rätt plats i utskottet för jordbruk och landsbygdens utveckling .
Innan kött , mjölk , bröd och andra produkter försäljs över disk kommer djurfoder och tillsatser att struktureras , blandas , mixas , skäras sönder och transporteras upprepade gånger .
Kampen bland djurfoderproducenterna för att uppnå största marknadsandel innebär , på samma sätt som inom livsmedelsproduktionen , många problem .
De negativa följderna känner vi till , de positiva vet vi mindre om .
Jag är fast övertygad om att hälsan för de europeiska konsumenterna i den ekologiska kedjan bäst kan skyddas genom att livsmedel och djurfoder produceras inom regionen och för regionen .
Men detta kräver ytterligare arbete .
Herr talman !
Får jag börja med att gratulera föredraganden , Graefe zu Baringdorf , för hans betänkande .
Det avspeglar åsikterna och oron hos alla EU-medborgare över frågor som rör livsmedelssäkerhet och livsmedelskvalitet .
Tidigare händelser under ett antal år har förvisso skapat en medvetenhet och farhågor om det verkliga hotet mot livsmedelssäkerhet och folkhälsa .
Den snabba insats som görs av detta parlament måste av alla medborgare anses som deras största garanti för framtiden för ni har lagt fast en dagordning om livsmedelskvalitet som medlemsstaterna måste rätta sig efter .
Men även på detta viktiga förvaltningsområde visar parlamentet sitt åtagande om subsidiaritet genom att uppmuntra medlemsstaterna att ta på sig sitt ansvar .
I Agenda 2000 har vi enligt min åsikt prioriterat politikområden som direkt berör medborgarna : livsmedelssäkerhet , vattenkvalitet , miljöskydd och utveckling av landsbygden .
Om vi fullföljer denna dagordning med engagemang och hårt arbete kommer de första åren av det nya millenniet att bli en milstolpe för genomförandet av en politik som är inriktad på människorna och som väldigt mycket speglar gemenskapens behov .
Jag välkomnar i synnerhet de föreslagna nya och strikta tillståndsförfarandena för tillsatser i djurfoder .
De som upptäcks bryta mot dessa måste behandlas strängt .
Jag gratulerar den nye kommissionären , Byrne , som ansvarar för livsmedelssäkerhet .
Han har en tung uppgift men har agerat snabbt och effektivt på kraven från denna kammare , liksom på konsumenternas oro .
Jag är särskilt glad att mitt eget land , Irland , ligger i frontlinjen med genomförandet av nya livsmedelsföreskrifter grundade på principen om spårbarhet .
Detta kommer att göra ön Irland till ett framstående centrum i framtiden när det gäller livsmedelsproduktion .
Herr talman , herr kommissionär !
Jag skulle också vilka gratulera föredraganden som har gjort ett utmärkt arbete och framför allt glädja mig åt den enhällighet som har rått på gruppnivå om detta ärende .
Det är således planerat att kommissionen skall byta ut de befintliga tillstånden mot tillstånd knutna till de ansvariga för saluföringen av tillsatserna genom en förordning och att dessa byten skall göras på samma gång i fråga om alla berörda tillsatser .
Vi måste återställa en sammanhållen rättslig ram .
Kommissionen föreslog att införa en rättslig grund från och med oktober 1999 i direktiv 70 / 524 / EEG för att ersätta tillstånden .
Vi måste emellertid se till att inte skapa snedvridningar av konkurrensen såsom Kindermann och Auroi påminde om .
Jag tror att vi också tydligt måste identifiera de genetiskt modifierade tillsatserna i djurfoder för att göra det möjligt för och garantera för slutkonsumenten att han kan välja GMO-fri mat eller mat baserad på GMO .
Konsumenten bör få behålla sin beslutsfrihet med full sakkännedom .
Detta förslag har ingen finansiell inverkan på gemenskapens budget , herr kommissionär .
Därför behöver vi för livsmedelssäkerheten en total öppenhet för producenterna och konsumenterna .
Jag är övertygad om att kommissionen kommer att kunna följa föredraganden som , vill vi påminna om , har uppnått enhällighet i utskottet för jordbruk och landsbygdsutveckling .
Herr talman !
Sedan BSE först dök upp har vi här i kammaren alltid sagt att djurfodret är en av de första och viktigaste beståndsdelarna för en säker produktion av livsmedel , för att skydda konsumenternas hälsa .
Därför gläder det oss att kommissionen lägger fram ett förslag om fodertillsatser .
Utskottet , som jag här talar för , nämligen utskottet för miljö , folkhälsa och konsumentskydd , beslutade i december - förutsatt att ordföranden i utskottet för jordbruk och landsbygdens utveckling i egenskap av föredragande skulle utarbeta ett sådant bra betänkande - att vi kan avstå från ett yttrande .
Trots detta vill jag säga ett par saker och ta ställning till några punkter .
Först kanske något om den rättsliga grunden .
Även om vi i parlamentet har en ny arbetsordning - och det mycket väl kan hända att det med den mycket ambitiöse ordföranden i utskottet för jordbruk allt oftare kan uppstå tvister mellan utskottet för jordbruk och utskottet för miljö när det gäller ansvarsområdet för lagstiftningen - är trots detta en sak helt klar för mig när det gäller sådana konflikter : Sammanhållningen i parlamentet är avgörande , och den rättsliga grunden i en fråga är avgörande för mig .
Därför - det måste jag säga er , herr Byrne - fördömer jag den rättsliga grund som valts .
Om den endast är en traditionell rättslig grund som övertagits från de tidigare direktiven , då är det fel att bibehålla den .
Amsterdamfördraget säger helt klart : När det gäller människors hälsa skall artikel 152 väljas som rättslig grund , och jag måste här säga till utskottet för rättsliga frågor och den inre marknaden i vår egen kammare : Det räcker helt enkelt inte att titta på kommissionens förslag och säga att det inte står någonting i det om hälsa och konsumentskydd , alltså handlar det inte heller om hälsa och konsumentskydd .
Därför kommer min grupp - som Kindermann redan sagt - i morgon att rösta för en ändring av den rättsliga grunden , och jag hoppas att de andra grupperna i kammaren också kommer att göra det .
Herr Byrne , jag ber er för öppenhetens och det goda samarbetets skull att anta och rösta för en ändring av den rättsliga grunden .
Om vi nämligen inte gör det , utan hörsammar utskottet för rättsliga frågor , skulle vi öppna dörren för manipulation .
Då tillåter vi nämligen kommissionen att välja den rättsliga grunden , så att politiken för folkhälsan helt enkelt inte nämns i texten , och då är det plötsligt fråga om artikel 37 .
Låt mig helt kort också säga något om de två andra punkterna : Beträffande genetiskt modifierade organismer i djurfoder får det inte vara så att man hänvisar till vertikal lagstiftning och säger att vi så småningom behöver en annan lagstiftning .
Men den har vi för närvarande inte !
Och så länge som vi inte har det , måste vi alltid när vi beslutar om lagstiftning också behandla genetiskt modifierade organismer , nämna dem särskilt och insistera på en märkning .
Det har föredraganden gjort , och det är ett bra tips .
Jag vill än en gång säga det som jag redan sagt många gånger : Ja , jag vill att kommissionen gör upp förslag till en positivlista .
Vi kommer säkert sedan att diskutera och behandla den kontroversiellt i denna kammare , men vi behöver åtminstone ha ett förslag till en positivlista för fodertillsatser .
Det är lika viktigt att vi har stränga hygieniska krav på produktionen av tillsatser och att det kontrolleras ordentligt i medlemsstaterna .
På båda områdena finns det fortfarande brister , och där har vi fortfarande mycket att göra .
Herr talman !
Jag vill gratulera föredraganden till hans betänkande .
Detta är en fråga som vi utan tvivel skall överväga på nytt vid flera tillfällen i framtiden .
Det som har hänt under de senaste åren har gjort oss uppmärksamma på de ofantliga problem som inte bara producenter av livsmedel utan även konsumenter kan vänta sig .
Vi måste hitta en balans mellan dem .
Vi måste lösa denna fråga eftersom det är viktigt att konsumenter återfår förtroendet för den mat de äter .
Ett sätt att uppnå detta är att införa total insyn när det gäller märkningen .
Genetiskt modifierade organismer ( GMO ) är den nya utmaningen för oss .
Detta är något som människor är mycket oroade över och helt med rätta och jag själv delar denna oro .
Men jag anser att vi inte skall tillåta vår oro över GMO överskugga vår oro över växtfrämjande ämnen i djurfoder eller antibiotika i foderblandningar .
I själva verket bör vi inte låta GMO skymma det faktum att kött- och benmjöl fortfarande ingår i djurfoder i många länder i Europa .
En faktor bakom denna utveckling som har nämnts i denna debatt är konkurrensen - konkurrens mellan medlemsstater om kostnaderna för livsmedelsproduktionen .
Detta är samtliga områden där vi måste säkerställa spelregler på samma nivå : livsmedel måste vara av samma standard i alla medlemsstater .
Vi har haft dioxinskräckupplevelsen , BSE och många andra problem .
Huvudproblemet är av ekonomisk art , nämligen vem bär kostnaden ?
Problemet är att kostnaden inte delas lika mellan konsumenten och producenten : producenten har tvingats bära alla kostnader .
Vi behöver en rättvis fördelning av de extra kostnader som uppstår .
Vi måste också se till att det livsmedel som importeras till Europeiska unionen håller samma standard som inom Europeiska unionen .
Om vi inte bibehåller dessa standarder för importerade livsmedel kommer vi att möta större svårigheter i framtiden . .
( EN ) Jag skulle först vilja tacka utskottet för jordbruk och landsbygdens utveckling och dess föredragande , utskottets ordförande , Graefe zu Baringdorf , för hans granskning av kommissionens förslag .
Kommissionens förslag är som några av er sagt ganska teknisk .
Ändå har den ganska enkla mål : att harmonisera förfarandena gällande tillstånd för fodertillsatser .
För närvarande skiljer sig handläggningen av tillstånd beroende på om ansökan lämnades före eller efter den 1 januari 1988 .
Syftet med kommissionens förslag är att harmonisera förfarandena för att kunna garantera att inga sådana skillnader finns .
Det föreslagna ändringsförslagets räckvidd är därför mycket begränsad .
Fem ändringsförslag har lagts fram av parlamentet .
Jag beklagar att kommissionen inte har möjlighet att godkänna dessa ändringsförslag trots det faktum att jag är helt medveten om uppfattningar och åtaganden hos parlamentet , utskottet för jordbruk och i synnerhet föredragande , Graefe zu Baringdorf , i dessa frågor .
Jag skall ta upp vart och ett av de enskilda ändringsförslagen separat .
I det första ändringsförslaget föreslås en ändring av den rättsliga grunden för förslaget och att ersätta artikel 37 med artikel 152 .
Jag vill endast påpeka att kommissionens förslag inte innehåller hänvisningar till hälso- eller konsumentskydd .
Den föreslagna ändringen är teknisk och kan inte tolkas ha som primärt syfte att skydda folkhälsan .
Jag konstaterar att parlamentets utskott för rättsliga frågor och den inre marknaden också godkänner att artikel 37 är den lämpliga rättsliga grunden .
Jag vill påminna parlamentet om att i artikel 152 är hälsoskyddet det primära målet .
Jag rekommenderar er de argument som anges i skrivelsen från utskottet för rättsliga frågor i vilken ståndpunkten fastslås med enligt min åsikt precision , tydlighet och med lovvärd kortfattad text .
Ändringsförslag 2 och 3 syftar mycket längre än kommissionens förslag eftersom syftet med dem är att införa ytterligare bestämmelser om genetiskt modifierade tillsatser .
Jag är den förste att gå med på att GMO är en mycket viktig fråga .
Jag godtar och erkänner också att ett antal initiativ för att aktualisera EU-lagstiftningen på området GMO krävs .
Detta tekniska ändringsförslag är emellertid inte det rätta instrumentet för att införa sådana initiativ .
Kommissionen anser att det är för tidigt att ändra de nuvarande fastslagna bestämmelserna i direktiv 70 / 524 om genetiskt modifierade tillsatser i detta skede .
I stället är det lämpligt att vänta på utvecklingen i förbindelse med den gemensamma ståndpunkten om ändringsförslag till direktiv 90 / 220 , vilken just nu är under den andra behandlingen i parlamentet .
Kommissionen planerar att gå mycket längre än vad som för närvarande föreslås av parlamentet i dess ändringar .
Jag kan även försäkra parlamentet att jag skall se till att de relevanta bestämmelserna i direktiv 90 / 220 innefattas i förslaget om en omarbetning av direktiv 70 / 524 som kommissionen föreslog i vitboken om livsmedelssäkerhet som skall läggas fram för parlamentet innan juli månad 2001 .
Jag kan också försäkra parlamentet att alla yttranden här i dag kommer att beaktas till fullo .
Ändringsförslag 4 och 5 kan inte heller godkännas för att de ger obefogat företräde till imitationsprodukter genom att bevilja tillstånd att omsättas till och med innan en ansökan om tillstånd har ingivits .
Kommissionen vidhåller att sådana ansökningar först skall bedömas i fråga om säkerhet och verkan innan tillstånd ges .
Jag kan bara be er igen att lägga på minnet den tekniska formen i kommissionens förslag och att avvakta det verkliga förslaget till ett nytt direktiv om fodertillsatser för att ta itu med större frågor .
Jag vill endast ta upp några av de specifika frågor som togs upp under debatten .
För det första , avseende synpunkter från herr Graefe zu Baringdorf , vill jag försäkra honom att vi kommer att ändra förfarandet för tillstånd till GMO tillsatser i tillsatsdirektivet 70 / 524 och inte i det nya foderdirektivet .
Detta är ett direktiv som mer specifikt behandlar råmaterial snarare än tillsatser .
Den text som parlamentet använde härrör från det direktiv som antogs 1998 .
Men den vertikala lagstiftningen i direktiv 90 / 220 om hur man bedömer miljörisker i samband med GMO har förändrats sedan dess och håller fortfarande på att förändras .
Det behandlas av parlamentet i en andra behandling .
Jag tror att vi bör vänta på det slutliga resultatet gällande direktiv 90 / 220 och i synnerhet , artikel 11 .
Man tog även upp frågan om detta förslag kunde skapa en risk för att monopol inrättades .
Kindermann och Auroi anspelade på detta .
Jag vill endast ta upp några punkter i den frågan .
För det första har detta ärende funnits i stöpsleven sedan 1993 , så det har faktiskt inte överrumplat några andra råvaruproducenter .
Varje sådan sökande kan i själva verket fortfarande lämna in en ansökan gällande sin speciella produkt .
Ja vill också understryka att kommissionen aldrig har godkänt någon ansökan om tillstånd att använda GMO i tillsatser .
Roth-Behrendt berörde frågan om lämplig rättsliga grund , om den borde vara artikel 37 eller artikel 152 .
Jag hänvisar återigen till vad jag sade tidigare om detta och försäkrar henne och kammaren att det skulle vara helt olämpligt för kommissionen att försöka försvara en åtgärd grundad på artikel 37 bara genom att i bestämmelsen undanta varje hänvisning till folkhälsa .
Detta är ett ärende som EG-domstolen behandlat vid minst två skilda tillfällen och den har fastlagt rättsliga kriterier för situationer som denna där lämpligheten hos den rättsliga grunden först måste prövas ordentligt när ny lagstiftning läggs fram .
Domstolens rättspraxis verkar helt klar med hänsyn till detta .
Som en generell kommentar till de här föreslagna ändringarna , särskilt med tanke på frågan om rättslig grund , skulle det vara olämpligt enligt min mening att ändra den rättsliga grunden till artikel 152 under dessa omständigheter då det är mycket troligt att det skulle komma i konflikt med de sakliga kriterier som domstolen lagt fast .
Fler av er - Nicholson i synnerhet - tog upp frågan om märkning .
I direktiv 70 / 524 förutses frågan om märkning av genetiskt modifierade tillsatser .
Det innehåller redan nu texten : " angivelse av särskilda karakteristiska egenskaper på grund av tillverkning av produkter " .
Således kommer denna fråga att tas upp .
Den formuleringen gjorde det möjligt för oss att ålägga sökanden att i märkningen ange det faktum att genmodifieringsteknik använts i produkten , sakinnehållet i ansökan . .
( DE ) Herr talman !
Tillåt mig ytterligare en fråga till kommissionären .
Först följande påpekande , kommissionär Byrne : Europaparlamentet har ingen initiativrätt när det gäller lagstiftningen .
Men när ni föreslår en ändring av ett direktiv eller en förordning tar vi oss rätten att titta på hela förordningen och inte bara på den del som ni valt ut .
Vi har dessutom i våra ändringsförslag begränsat oss till en formell tillnärmning till andra direktiv .
De innehållsliga frågorna har vi till och med avstått från .
De går till exempel inte in på antibiotika .
Därför handlar det bara om tillnärmning av de rättsliga bestämmelserna i de enskilda direktiven .
Min fråga , kommissionär Byrne : Vid FN : s konferens i Montreal har man just genomdrivit att det i det internationella handelsutbytet måste finnas en märkning av genetiskt modifierade organismer .
Tror ni verkligen , att parlamentet - när vi nu har denna möjlighet - kan tillåta att denna märkning inte genomdrivs inom Europeiska unionen för fodertillsatser ?
Kommissionär Byrne , ni är på väg mot en kraftmätning med parlamentet .
Vi har förhandlat om lagen om utsäde i två år .
Jag ser fram emot våra gemensamma diskussioner . .
( EN ) Jag vill bara understryka att inga genetiskt modifierade organismer har godkänts enligt detta direktiv ; det gäller enbart för tillsatser .
Jag vill också säga beträffande frågorna om märkning att detta är en komplicerad fråga .
Man håller på att granska detta och skall undersökas på ett allsidigt sätt , särskilt i direktiv 90 / 220 .
Denna fråga behandlas just nu av parlamentet och det kommer att bli andra direktiv rörande denna fråga som också kommer att ha artikel 152 som rättslig grund , vilket ger parlamentet fullständig behörighet i fråga om medbeslutande .
Jag vill försäkra herr Graefe zu Baringdorf att det inte alls är min avsikt att få någon sammandrabbning eller styrketest med parlamentet i denna fråga .
Min avsikt är som den alltid har varit att samarbeta med parlamentet , att se till att de resultat som vi uppnår är de absolut bästa resultaten .
Det bästa sättet att lösa denna fråga är för närvarande genom att lägga fram lagstiftningsförslag för parlamentet , liksom lagstiftningen under utarbetande , snarare än i detta tekniska dokument och under förhållanden där man kanske inte helt har tagit hänsyn till de frågor som läggs fram och som skall diskuteras inom ramen för direktiv 90 / 220 .
Det är bäst att avvakta den debatten som enligt vad jag hört skall ske ganska snart .
Alla dessa frågor skall tas upp i det lagstiftningsarbetet .
Tack , herr kommissionär .
Parlamentet noterar era anmärkningar .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.30 .
 
Skrapie Nästa punkt på föredragningslistan är betänkande ( A5-0023 / 2000 ) av Böge för utskottet för jordbruk och landsbygdsutveckling om förslaget till Europaparlamentets och rådets direktiv om ändring av rådets direktiv 91 / 68 / EEG i fråga om skrapie ( KOM ( 1998 ) 623 - C4-0026 / 1999 - 1998 / 0324 ( COD ) ) .
Herr talman , herr kommissionär , kära kolleger !
Det har alltid hört till egendomligheterna och de gåtor som hittills inte lösts när det gäller bearbetningen av BSE-affären att vi hittills inte haft några gemenskapsregler för bekämpning av skrapie hos får .
Därför hörsammar kommissionen absolut med sina förslag att ändra direktiv 91 / 68 och stryka hänvisningen till skrapie - även med tanke på kollegan Roth-Behrendts betänkande som också skall diskuteras här om förebyggande och bekämpning av TSE-infektioner generellt - också parlamentets krav , som bygger på den efterbearbetning som gjorts av det tillfälliga utskottet för uppföljning av rekommendationerna beträffande BSE .
Vi välkomnar detta eftertryckligen .
Här vill jag emellertid också tillfoga att det inte hade krävts några nya forskningsrön som gav belägg för att en experimentell infektion av får genom utfodring med BSE-material leder till kliniska manifestationer , som inte skiljer sig från kännetecknen på skrapie-sjukdom .
Dessa nya rön hade inte krävts , eftersom man redan från början baserat sig på den alltmer etablerade teorin , att BSE mycket väl måste ha något att göra med skrapie .
Därför har vi har vi blivit litet försenade .
Jag kan alltså absolut rösta för kommissionens förslag vad gäller skrapie .
Men jag vill också tillfoga , att detta bara är meningsfullt om vi i den kommande nya TSE-förordningen strikt gör en förnuftig symbios av konsumentskyddet och förslagens genomförbarhet .
Därför kommer det också i den kommande debatten om TSE-förslaget - hela tiden också med beaktande av skrapie - an på att vi egentligen konsekvent tar hänsyn till sex - sju punkter .
När vi talar om TSE-förordningen hör det också hit , herr kommissionär , att det klargörs att vi beträffande produkter som är undantagna från denna förordning , exempelvis kosmetika , läkemedel och även kött- och benmjöl , mycket snabbt kommer fram till särskilda förslag på grundval av motsvarande rättslig grund , artikel 152 .
Det insisterar vi på .
För mig hör det också hit att de helt grundläggande kärnbestämmelserna i detta förslag till förordning inte får återfinnas i bilagan , utan de hör hemma i förslaget till förordning som sådant , eftersom vi som parlamentet här vill och kommer att ta del i ansvaret .
Det är också så att i fråga om bekämpningen hör problemet med undantag av hela hjordar i samband med skrapie eller BSE-angrepp fortfarande till föredragningslistan , och likaså frågan om avgränsning av geografiska områden .
Även om jag välkomnar att skrapie-bekämpningen tas upp i TSE-förordningen anser jag fortfarande att kommissionens förslag med tanke på bekämpning av skrapie inte är tillräckligt konsekventa .
Därför kommer jag att lämna in förslag i samband med Roth-Behrendts betänkande , även för utskottet för jordbruk och landsbygdens utveckling , som kommer att leda till en skärpning .
Dessutom vill jag beröra ytterligare två punkter : Vi välkomnar eftertryckligen principen med regionalisering av medlemsstaternas statusklasser med tanke på skrapie- eller TSE-angrepp .
Även här har kommissionen alltmer hörsammat parlamentets arbeten och krav .
När vi avslutningsvis talar om den kommande användningen av tester , måste vi naturligtvis veta att vi ännu inte kommit så långt att testerna kan utvärderas generellt .
Men de tester som man i dag förfogar över är ju absolut lämpade , visserligen inte att för varje enstaka djur garantera konsumenterna någon hälsopolitisk säkerhet , men när det gäller att tala om huruvida en region kan överflyttas från en negativ status till ett mer gynnsamt läge i fråga om bekämpning av djursjukdomar kan den epidemiologiska granskningen av situationen i en region , genom lämpliga stickprov i slakthuset då man använder sig av sådana tester , visa på en klok väg även i den politiska och vetenskapliga debatten , där vi iakttar förebyggande konsumentskydd och i grund och botten , genom att använda sådana tester , också kan lösa konflikter på en ordentlig grundval bättre än vad som tidigare varit möjligt .
Jag ber er , herr kommissionär , att redan nu ta med er dessa reflexioner så att säga på väg till betänkandet om skrapie och till det generella bekämpningsbetänkandet om TSE , och ställa in er på att vi kommer att fordra dessa punkter av er .
( Applåder ) Herr talman !
Under tidens gång har följande situation uppstått : En fråga har nu under flera år vidareutvecklats i de mest skilda varianter .
Många av oss här i kammaren har i många år - vare sig de ville eller inte - i stor utsträckning inte ägnat sig åt något annat än konsekvenserna av BSE-skandalen , ända fram till de sista varianterna .
Det är i dag fortfarande ett ämne .
Därför är det ju heller inte underligt att Böge och jag talar om det , och att Graefe zu Baringdorf också just har nämnt det i sitt betänkande .
Det är ju samma agerande personer .
Det är säkerligen - även om orsaken var otrevlig - inte den sämsta erfarenhet som detta parlament gjort .
Min uppgift som föredragande av yttrandet från utskottet för miljö , folkhälsa och konsumentpolitik är mycket enkel .
Jag kan hålla med föredraganden och säga att utskottet har bett och krävt av utskottet för jordbruk och landsbygdens utveckling att man skall rösta för kommissionens förslag .
Därigenom har jag vunnit mycket tid , som jag ibland gärna vill använda för andra saker , och som jag nu litet grand i förväg också vill utnyttja , som Böge redan har gjort .
Mitt betänkande om TSE har kammaren ännu inte fått .
Vi var till att börja med litet obeslutsamma , även om vi beklagar det .
Men jag har kommit fram till att det egentligen är en ganska bra " timing " .
Det är egentligen riktigt bra att vi med ledning av denna debatt också redan nu kan ge kommissionen ett par saker att tänka över , herr Byrne .
Efter att vi kanske tidigare , när det gällde Graefe zu Baringdorfs betänkande , inte behandlade varandra så positivt och säkert inte heller kommer att närma oss varandra särskilt mycket , så kan det ju hända att det i fråga om detta betänkande blir litet annorlunda .
Låt mig redan nu säga att den del av det komplexa betänkande , som Böge har behandlat - för övrigt är det en bra form av samarbete mellan två utskott , att man låter det ena utskottet vara ansvarigt , medan det andra avger ett yttrande , och tvärtom , vilket kanske kan vara ett exempel för framtiden - är relativt enkelt .
Svårare blir det när vi kommer att titta på TSE-förslaget , herr Byrne .
När vi då ställer direkta frågor , kommer de frågor upp som Böge redan har berört .
Då kommer frågan - och den kommer jag att tvingas ställa till er och även till kommissionens företrädare i utskottet - hur det kommer att se ut med BSE-statusen i medlemsländerna och i tredje land .
Hur kommer BSE-statusen faktiskt att definieras ?
Kommer ni eventuellt också vara beredda att använda en BSE-test när det gäller BSE-statusen ?
Och sedan min ständiga fråga till er , herr Byrne , som ni ju säkert redan känner igen och som inte heller överraskar er : Hur är det nu med BSE-testen ?
När kommer ni att göra den obligatorisk ?
Kanske gör ni det rent av innan detta parlament diskuterar TSE-betänkandet .
Jag vill inte förhala det , men det skulle ju så att säga vara en fin gest , om ni kunde säga : Och här har ni nu lagstiftningsförslaget om BSE-testerna !
Jag vet att jag plågar er med detta , herr Byrne , men ibland måste det göras .
Jag vill eftertryckligen säga - och detta också efter Graefe zu Baringdorfs betänkande , som ju är starkt förknippat med hela idén - att djurfoder , djurhållning och djurproduktion måste vara sådana att de för det första är anpassade efter arterna , och för det andra måste de framför allt vara sådana att människorna inte skadas eller utsätts för risker .
Det får ändå inte vara så att ni undantar kosmetika , farmaceutika och andra produkter med motiveringen att det inte kan uppstå några skador eller att det inte är farligt .
Det är med säkerhet för kort , för knappt och för litet sagt .
Ni har tur eftersom detta i Böges betänkande behandlas i periferin .
Men beträffande mitt betänkande kommer ni att få det problemet att ni måste rättfärdiga er litet bättre , och ni kommer att få litet mer problem med det .
Avslutningsvis också ett kort påpekande , herr Byrne .
Vi har en ny kommission .
Om vi i framtiden kommer att vara införstådda med denna kommissions och med kommissionsordförandens arbete , det får tiden utvisa .
En sak kommer vi säkert inte att kunna överse med , och det kan ni som jurist och politiker nog förstå : Det får inte vara så att det som verkligen är det viktiga , regleras i bilagor .
Det hör till lagstiftningstexten .
Om jag vore kommissionär , skulle jag kanske också göra på så vis , eftersom jag på ett enkelt sätt kan ändra en bilaga med hjälp av kommittéförfarandet , och jag inte alltid måste samarbeta med detta parlament , som behöver så lång tid på sig och också är så svårt att samarbeta med .
Men ni måste förstå att vi inte kan ha överseende med detta .
Det betyder att så snart jag kan påverka , så hämtar jag ut allt ur bilagorna och sätter in det i lagstiftningstexten .
Det är alltså bäst att ni gör det redan från början !
( Applåder ) Herr talman !
Herr kommissionär !
Mina damer och herrar !
Jag vill i dag erinra om hur vår livsmedelskedja är sammansatt och hur viktigt det är att denna kedja ger människorna säkra och hälsosamma livsmedel .
Produktionen måste utan undantag vara fri från tvivelaktiga och riskabla mellan- och slutprodukter .
Under de senaste åren har dessa grundprinciper på grund av slarv eller girighet ignorerats inom djurhållning , djurutfodring och också ofta även när det gäller djurhälsovillkor .
Europaparlamentet har redan intagit en klar hållning i fråga om BSE , och jag anser att detta borde vara fallet i fråga om alla djursjukdomar .
Vi får inte låta någonting skada livsmedelssäkerheten , ty det handlar i sista hand om vår hälsa .
Kommissionens förslag omfattar inte bara transport och avyttring av får och getter , utan även gemenskapsbestämmelser för bekämpning av skrapie .
Detta är desto viktigare som vi ännu inte har något entydigt besked om att det inte finns något sammanhang mellan BSE och skrapie .
Det köps djur i hela Europa som transporteras över kontinenten .
Epidemier som sprids på grund av att ett sjukt djur förs in kan få oerhörda följder för jordbrukarna .
Och jag vill påpeka att det för första gången i historien uppträtt ett skrapie-fall också i Österrike .
Skrapie är en särskilt lömsk sjukdom , eftersom sjukdomsalstrarna kan ligga aktiva i dammet i flera år , och åter tas upp via fodret .
Sjukdomen leder alltid till döden .
Eftersom det inte heller är möjligt att vaccinera mot den , kan en jordbrukare bara skydda sig genom att inte köpa några djur från länder med skrapie-fall .
Även om skrapie inte kan överföras till människor , så är sambandet med BSE - som redan sagts - fortfarande oklart .
Man får inte skapa några risker för konsumenten , detta ligger mig som jordbrukare mycket varmt om hjärtat .
Jag förespråkar att man vidtar förebyggande åtgärder , som börjar med ett artanpassat djurfoder , i stället för åtgärder för att bekämpa en epidemi som redan brutit ut .
Jag välkomnar därför kommissionens initiativ att skapa en ny rättslig grund för bekämpningen av skrapie .
( Applåder ) Herr talman , ärade kommissionär !
Böges betänkande om åtgärder för bekämpning av TSE-sjukdomar hör till de frågor som bygger på de förslag som framförts av parlamentets tillfälliga BSE-utskott .
Böge har gjort ett betydelsefullt arbete i detta utskott och det är en lättnad att se att det är han som fått i uppdrag att följa upp BSE-utskottets arbete i utskottet för jordbruk och landsbygdens utveckling .
Han har erfarenhet .
Jag hade gärna kommit med ett anförande i den diskussionen om man samtidigt hade diskuterat den andra delen av kommissionens förslag .
Jag tycker inte det är ändamålsenligt att vi delvis måste föra samma diskussion igen då vi får Roth-Behrendts betänkande från utskottet för miljö , folkhälsa och konsumentskydd till kammaren .
I föregående inlägg konstaterade Schierhuber att skrapie är en mycket förrädisk sjukdom .
Det stämmer .
För mig som finländare , som har arbetat nära jordbruket i frågor som rör djurens hälsa och transport av djur , är det viktigast att de länder där TSE-sjukdomar inte alls förekommer också i fortsättningen garanteras rätten att i tillräcklig grad granska transporter av levande djur .
Möjligheten att vid behov granska djuren ytterligare inom dessa områden är inte någon konstgjord protektionism eller någon begränsning av den fria rörligheten när orsaken är välmotiverad .
Granskningarna måste ses som rättvisa och kostnadseffektiva handlingar med vilka man främjar djurens välbefinnande och förhindrar att nya kostnader uppstår för EU .
För Europeiska liberala , demokratiska reformistiska partiets grupps del kan vi godkänna kommissionens förslag i den mån det gäller Böges betänkande , men i behandlingen av nästa betänkande av Roth-Behrendt måste vi på nytt återgå till situationen i de länder , där TSE-sjukdomar inte förekommer .
Herr talman !
Även jag vill gratulera föredraganden .
Det finns inga tvivel om att Böge och föredraganden för utskottet för miljö , folkhälsa och konsumentfrågor nu är fantastiska experter på detta område .
Det är mycket bra att de fortsätter att bevaka denna fråga på parlamentets vägnar eftersom den är ytterst viktig .
Oavsett de många andra angelägna frågor vi har har BSE gett oss ett fruktansvärt arv som måste hanteras och lösas .
Det är helt klart att förekomsten av skrapie hos får har varit en bidragande orsak till hela problemet .
Jag är positiv till den rättsliga grund som läggs fast och till det samlade sättet kommer de nya bestämmelserna hoppas jag att kunna lösa denna situation .
Vi måste kunna garantera att ingenting kan införas i livsmedelskedjan eller i djurfoderblandningar så att vi inte låter det som vi tidigare varit med hända på nytt i framtiden .
Ingen skulle vilja se att det som hände för bönder med BSE någonsin kunde hända igen .
Vi måste tillämpa de mest strikta bestämmelser och vi måste få dem att fungera .
Det är ytterst viktigt både för producenten och konsumenten att vi återställer förtroendet och det enda sättet vi kan göra det på är genom att ytterst noggrant ta itu med problemet och lösa det .
BSE har verkligen inte försvunnit .
Man kan hitta det i olika länder .
Jag vill inte peka på något speciellt land men många länder står nu inför liknande problem som dem vi hade i Förenade kungariket .
Den kommer att finnas kvar under ytterligare någon tid .
Vi måste se till att hela systemet med spårbarhet och möjligheten att följa djuret från födsel till slakt och rakt genom hela livsmedelskedjan blir en del av den förtroendeskapande mekanismen .
Om vi inte kan uppnå det kommer vi att få ofantliga problem i framtiden .
Till sist , eftersom jag själv har jordbruksbakgrund har jag under en lång tid absolut trott att om vi hade utfodrat djuren med rätt foder och om djurfodret hade framställts av rätta blandningar skulle vi aldrig haft BSE för det första .
Det handlade aldrig om bondens ansvar utan det var producenterna av foderblandningar som orsakade detta problem och vi måste försäkra oss om att det aldrig händer igen . .
( EN ) Herr talman !
Jag är glad att jag fått detta tillfälle att diskutera en fråga där det finns ett gott samarbete mellan parlamentet och kommissionen , nämligen att bekämpa TSE .
Jag vill också tacka herr Böge för hans arbete i denna fråga .
Betydande framsteg har gjorts om vårt förslag till Europaparlamentets och rådets förordning om skydd mot och kontroll av TSE enligt artikel 152 i fördraget .
Detta förslag innehåller alla TSE-risker i alla djur och i alla faser i produktionskedjan .
Jag är här i dag för att lyssna på era synpunkter på det första steget i denna process för att införa en verkligt omfattande gemenskapssystem för att kontrollera dessa sjukdomar .
I det aktuella förslaget har jag föreslagit att man skall stryka alla nu gällande gemenskapsbestämmelser om skrapie hos får och getter och att införliva dem i ramförslaget om en förordning .
Närmare bestämmelser skulle då läggas fram i det ramförslaget .
Jag har informerats om att ni är positiva till detta initiativ , vilket verkar vara fallet enligt era bidrag denna eftermiddag , att utforma en enda text .
Jag ser fram emot att diskutera varje ytterligare förbättring ni önskar föreslå enligt ramförslaget till lagstiftning , särskilt efter den hänvisning som Roth-Behrendt gjorde till sitt eget betänkande och ståndpunkt i denna fråga .
Jag ser fram emot att få det dokumentet som kommer att beaktas vid alla ytterligare överväganden med hänsyn till denna fråga .
Till sist vill jag framföra detta rörande synpunkten att föra in lagstiftningen i bilagor och synpunkten att vi måste uppnå en effektiv balans mellan parlamentets rätt att lämna sina synpunkter och samtidigt vårt krav om snabba resolutioner , snabb lagstiftning och snabba ändringar till gällande lagstiftning .
Under de månader jag har varit kommissionär och sett hur lagstiftningsarbetet fungerar i hela systemet inser jag att det krävs mycket arbete på detta område så att vi alla kan uppnå det vi strävar efter , det vill säga överföring av politik till lagstiftning .
Tack , herr kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.30 .
 
Gemenskapsåtgärder på vattenpolitikens område Nästa punkt på föredragningslistan är andrabehandlingsrekommendation ( A5-0027 / 2000 ) om rådets gemensamma ståndpunkt ( 9085 / 3 / 1999 - C5-0209 / 1999 - 1997 / 0067 ( COD ) ) inför antagandet av Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder på vattenpolitikens område ) .
( Föredragande : Marie-Noëlle Lienemann ) . .
( FR ) Herr talman , mina damer och herrar kommissionärer , kära kolleger !
Vattenfrågan kommer att vara en av de stora miljö- och världsfrågorna under det tjugoförsta århundradet .
Om det så handlar om klimatförändringar , världsövergripande resurser , kvaliteten i våra floder och kvaliteten i våra underjordiska vatten , vet vi att de stora utmaningarna medför risker för vår gemensamma framtid .
Antingen kommer vi att kunna återställa en vattenkvalitet som motsvarar jordens ekosystem eller så kommer vi att få se en hel rad störningar som hotar utvecklingen i vissa områden och som hotar invånarnas livsvillkor i andra områden , och i grund och botten till och med den globala jämvikten .
Som bevis använder jag en utmärkt rapport som vår kollega Mario Soares har upprättat i de internationella instanserna om havens och oceanernas tillstånd .
När vi talade om klimatförändringar hänvisade vi med rätta till växthuseffekten och atmosfärens tillstånd .
Men vi vet också att försämringen av oceanerna i hög grad kommer att destabilisera stora delar av vår jord .
Europa bör lämpligen vara så att säga exemplariskt i sina metoder både för att det bör främja en viss modell för utveckling och för att det själv står inför allvarliga problem med föroreningar och vattenförsämring , vare sig det handlar om underjordiska vatten , ytvatten eller hav .
EU har för övrigt undertecknat internationella konventioner .
Jag tänker särskilt på Ospar-konventionen ( International Commission for the Protection of the North East Atlantic ) genom vilken EU har gjort åtaganden .
EU sade " om några år bör vi ha stoppat utsläppen av föroreningar , vi bör ha upphört med att öka föroreningarna och bör till och med närma oss nollstrecket i fråga om giftiga eller farliga ämnen " .
EU undertecknar således de internationella avtalen , därefter följer ett direktiv samt konkreta politiska åtgärder ute i terrängen och då meddelar EU att de fastställda målen inte kommer att kunna uppnås eller också skjuts de upp till sådant datum att själva trovärdigheten i undertecknandet av de internationella avtalen ifrågasätts .
När Europaparlamentet tog upp debatten om ramdirektivet om vattenpolitik ansträngde parlamentet sig därför redan vid första behandlingen att kräva en sammanhållning mellan ramdirektivet och de internationella målen samt i synnerhet , när det gäller respekten för Ospar , en konvergens som är effektiv och konkret samt stimulerar oss till åtgärder .
EU : s vattenpolitik utgår inte från ingenting .
Många direktiv har antagits och kommissionens vilja är för övrigt att lyckas med att göra dem läsbarare , mer överensstämmande sinsemellan samt förse dem med tydligare mål .
Det är således en rationell vilja som har lett till genomförandet av detta ramdirektiv .
Men parlamentet insisterade vid första behandlingen på att det aktuella direktivet inte bara skall överensstämma med våra åtaganden - typ Ospar - utan göra det möjligt för oss att vända på utvecklingen .
För , trots de många direktiven och trots de upprepade förklaringarna om den ansträngning som bör göras i fråga om vattenskydd , när vi ser på miljösituationen i Europa , kan vi notera att målsättningarna inte har uppfyllts .
I många fall har situationen förvärrats och vi kan således inte nöja oss med en ansträngning att rationalisera texterna Vi bör sätta upp mål i nivå med de utmaningar som vi har framför oss , och vi har inte mycket tid på oss , för om vi tar för långa frister , såsom kommissionen hade föreslagit , kommer vi inte bara att få ett trovärdighetsproblem hos allmänheten , utan vi vet mycket väl att ansträngningarna kommer att skjutas upp till senare , därefter kommer de att skjutas upp på nytt och således vet man att man inte kommer att nå de uppsatta målen .
Jag trycker på denna punkt , för vi får inte vänta oss för hundrade gången att katastrofer rapporteras varje dag i våra tidningar för att säga " jaså !
EU har inte gjort det , jaså !
EU borde ha ... " och då skynda oss att låtsas lösa de problem som man inte ville ta itu med i rättan tid .
Exemplet för närvarande med Donau och den förorening som sker i Rumänien visar mycket tydligt att om vi inte inför en ny ekonomisk utvecklingsmetod , tydliga krav , kontroller och vidtar exakta åtgärder för våra floders tillstånd , vet vi att denna typ av olyckshändelse inte bara kommer att upprepas utan kommer att mångfaldigas med tiden .
Vi vet också att om vi inte gör någonting kommer utvecklingen av jordbruket att fortsätta att skapa stor obalans .
Floderna i Bretagne i mitt eget land är redan nu i en situation av total eutrofiering och det skadar turismen .
Herr talman , jag skulle bara vilja avsluta med att säga att det som står på spel är fullt ut klargjort i den andra behandlingen .
Vill vi , ja eller nej , ha normer som är förenliga med Ospar , det vill säga närma oss noll när det gäller farliga ämnen ?
Vill vi förkorta de frister som rådet har föreslagit för detta direktiv ?
Vill vi ha en prispolitik som ger möjlighet åt samtliga offentliga och privata aktörer att minska föroreningarna , att verka för föroreningsminskningar och spara vårt vatten ?
Vill vi seriöst uppfylla folkens önskningar ?
De flesta ändringsförslag som godkändes av utskottet för miljö , folkhälsa och konsumentfrågor uppfyller denna målsättning , jag hoppas att de kommer att få kammarens stöd .
Herr talman , mina damer och herrar !
Lienemann har ju nyss redan på ett drastiskt sätt förklarat hur viktigt det är för oss med vatten och luft , framför allt just som grundval för livet för oss människor .
Förutom vattenkvaliteten handlar det också om vattenmängden , ty det finns inte heller tillräckligt med vatten överallt i Europa , framför allt inte i de mycket torra områdena .
Jag beklagar att jag för ögonblicket inte kan se kommissionär Wallström här , som egentligen är ansvarig , ty det är hur som helst ett synnerligen viktigt direktiv , som kommissionen har arbetat mycket länge på , och den vattenskyddslagstiftning som vi i dag diskuterar i den andra behandlingen berör alla medborgare i Europeiska unionen , men också alla människor i kandidatländerna , som ju måste uppfylla EU : s lagstiftning när de ansluter sig .
Vi har arbetat i tio år med denna fråga , och den omfattande ansatsen har blivit möjlig först genom en utfrågning som initierades och genomfördes av utskottet för miljö , folkhälsa och konsumentfrågor .
Från den tidpunkten fram till den andra behandlingen i dag har många deltagare i Europaparlamentet , kommissionen och ministerrådet arbetat hårt med den .
De 243 ändringsförslagen i utskottet för miljö har vi reducerat till 77 , men nu har ytterligare 30 tillkommit .
Ni ser att det finns många frågor , och frågorna är av olika art .
Somliga vill ha en skärpning , andra en precisering , många är nationellt präglade .
Också i min grupp , Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokrater , har vi naturligtvis haft olika synpunkter .
Vi strävar efter realistiska mål och genomförbara lösningar .
I den andan betyder de ändringsförslag som jag och några kolleger har lagt fram från gruppens sida absolut en förbättring av de krav som föreskrivits i den gemensamma ståndpunkten .
Vissa ändringsförslag som vi stöder skall stärka Europaparlamentets förhandlingsposition i den kommande förlikningen med ministerrådet .
Vi säger klart nej till alla orealistiska krav , som skulle göra Europaparlamentet ovederhäftigt .
Hit hör för mig nollkravet , dvs. kravet på nollutsläpp fram till år 2020 .
Det skulle innebära slutet på all jordbruksverksamhet och mycket av industriverksamheten .
Här vill jag än en gång särskilt betona att med de befintliga nationella och europeiska lagarna till skydd för vattnet , hur ofullständiga de än varit och hur litet de än beaktats i medlemsländerna , har vi trots detta redan gjort avsevärda framsteg .
Jag vill bara erinra om att vi i dag åter har lax i Rhen , vilket för 20 år sedan fortfarande hade varit otänkbart , och att det denna vår skall sättas ut lax till och med i Elbe , som varit särskilt förorenad .
Det betyder ej att vi inte även i fortsättningen måste göra väldiga ansträngningar för att fortsätta att förbättra skyddet för vattnet och bibehålla den goda vatten- och grundvattenkvalitet som ännu finns , vilket naturligtvis utan tvivel också kommer att vara förbundet med avsevärda kostnader .
Många farhågor har just under de senaste dagarna yttrats från jordbrukets sida .
Också jordbruk kan bara bedrivas om det finns tillräckligt med friskt vatten till förfogande .
Med den linje som vår grupp följt för förhandlingarna med ministerrådet kommer man också att uppnå en bra lösning för jordbruket .
Jag bedömer att ledamöterna och allmänheten i detta svåra och delvis mycket tekniska ämne har vilseletts med falska argument från båda sidor .
Jag tackar därför i synnerhet mina kolleger i gruppen , som har bidragit med kompromisser .
Jag tackar särskilt vår föredragande Lienemann för hennes enorma arbete och hennes samarbetsvilliga hållning , även om det fortfarande finns olika uppfattningar på vissa punkter .
Men jag tackar också företrädarna för kommissionen , som hela tiden har bistått oss med råd och experthjälp .
Om företrädarna för ministerrådet intar en liknande konstruktiv hållning , betvivlar jag inte att vi alla gemensamt kommer att uppnå en ännu bättre lösning för vattenskyddet i Europa under förlikningen .
Herr talman !
Jag vill börja med att gratulera Lienemann till det utmärkta arbete som hon har lagt fram och till hennes ansträngningar för att närma våra skilda ståndpunkter i vattenfrågan .
Ramdirektivet om vatten är ett nödvändigt initiativ .
Om man däremot utgår från att tanken på solidaritet är en reell tanke för processen med det europeiska bygget , är det nödvändigt att man i direktivet tar hänsyn till att vattenresurserna betraktas som en faktor för den sociala sammanhållningen .
Vatten - det är det ingen som betvivlar - är en resurs av allmänt intresse .
Hanteringen av vattenresurserna förutsätter dock politiska lösningar , när det gäller Spanien och andra länder söderut med ett oregelbundet klimat , för att rationalisera förbrukningen samt andra åtgärder för solidaritet .
Vi anser att man i detta direktiv bör förespråka en användning av vattnet som gör det möjligt att åtgärda den territoriella obalansen och därför ber jag att ni stödjer ändringsförslag 95 , som har lagts fram av vår grupp .
Vi vill säkerställa att artikel 1 i direktivet främjar en hållbar , effektiv , rättvis och solidarisk användning av vattnet .
Jag vill nu göra en kort genomgång av de viktigaste punkterna där den spanska socialistiska delegationens uppfattning skiljer sig från de åsikter som försvaras här .
Det gäller överföring av vatten mellan magasin .
Vi anser att det vore bättre att ett framtida ramdirektiv inte innebar att möjligheten att genomföra dessa är föremål för gemenskapens övervakning .
Vi anser med tanke på den spanska statens säregna vattensituation , där överföring sker av strukturell natur , att det bör vara landets myndigheter som beslutar om det egna landets resurser , ett beslut som naturligtvis alltid skall grunda sig på kriterier med sammanhållning och en rationell användning av vattnet som målsättning .
Vad beträffar en av de mest omdiskuterade frågorna i vår debatt , nämligen prissättningen , har de spanska socialdemokraterna länge försvarat tanken att direktivet , alltifrån respekten för principen om att " förorenaren betalar " , skall förespråka en policy med rimliga priser på samtliga förbrukningsnivåer .
Det är uppenbart att en policy med ett fullständigt återvinnande av vattenkostnaderna inte skulle få samma effekt i Spanien som i länderna i centrala och norra Europa .
För spanjorerna skulle det innebära att kostnaderna för vattnet ökade för användningen på olika områden , just på grund av de bristande vattenresurserna och för att miljökostnaderna måste inbegripas inom ramen för det som direktivet fastställer .
Därför har vi alltid försvarat ett progressivt system för återvinning av kostnaderna , ett system där man har de sociala , miljömässiga och ekonomiska effekterna i åtanke , ett system vars tillämpning anpassas till de olika geografiska och klimatmässiga omständigheterna .
Vi vill bygga ett Europa med en hållbar och hälsosam omgivning .
Men ett miljövänligt Europa kan under inga omständigheter byggas i olika hastigheter , utan det bör byggas på en solidarisk grund .
Herr talman !
Den ekologiska katastrofen i Donau påminner oss om hur nära alla länder i Europa hör samman och hur viktigt vattnet är för oss alla .
Utflödet från kemiska fabriker i min egen valkrets i nordvästra England kommer till slut att hamna på stränderna på Europas fastland .
Detta klargör de samband som binder oss tillsammans .
Detta ramdirektiv är avsett att måla upp en bred skiss för vår politik under de kommande decennierna och det har funnits mycket panik rörande detaljerna .
Det är viktigt för oss att komma ihåg att detta är rambestämmelser .
Denna skiss är i själva verket mycket generell .
Det är lätt för enskilda länder , för enskilda industrisektorer att undkomma de effekter som har målats upp för oss under de senaste dagarna .
Det finns många möjligheter att komma undan .
I verkligheten kommer närmare bestämmelser i denna lagstiftning att fastläggas i dotterdirektiv för månader och år framöver .
Då är rätta tiden att diskutera några av dessa detaljproblem .
De breda principerna är verkligen sådana som vi borde kunna godkänna - de breda principerna att vi vill minska spridning av riskavfall till grundvattnet , de breda principerna att vi bör inrikta oss på att se till att de kemikalier som vi alla behöver i samhället under alla förhållanden inte bör kunna läcka ut i våra vattensystem .
Det finns en kemisk fabrik i nordvästra delen som skrev till mig för att säga att vi måste rösta emot denna lagstiftning .
Jag måste fråga dem vad det är för kemikalier som de släpper ut i vattensystemet just nu , och varför de inte meddelar alla som bor i det området exakt vad de håller på med .
Detta är något som de helst vill undvika att göra .
Principen gäller även vattenhushållning .
Den grundläggande insikten som många av oss nu delar är att vi måste införa miljöbeskattning för att uppmuntra till bevarande av resurser , att använda morot och sticka för att få alla att använda våra tillgångar på bästa sätt så att vi inte bidrar till ökad miljöförstöring eller en minskning av en så värdefull resurs som vatten .
Jag vill kommentera den politiska positionen här .
Den gemensamma ståndpunkten har gjort den ståndpunkt som intogs av parlamentets svagare vid första behandlingen .
Några icke-statliga organisationer skulle säga att direktivet i sin nuvarande utformning är sämre än värdelös .
Det är ett steg tillbaka .
Detta är en möjlighet för oss att förbättra situationen .
Vi måste vara i stånd att inleda ett medlingsförfarande .
Vi har sett omröstning efter omröstning förloras .
Åtgärd efter åtgärd har kommit från utskottet för miljö , folkhälsa och konsumentfrågor .
Vi har misslyckats med att skapa kvalificerad majoritet .
Våra försök att förbättra Europas miljö har misslyckats .
Vi måste försöka få till stånd ett medlingsförfarande .
Vi behöver i slutet av dagen kunna vara säkra på att vi slutligen får en klok och avvägd politik av verkliga förbättringar till rimliga kostnader .
Herr talman , kolleger !
Redan för nästan trettio år sedan försökte Europeiska kommissionen slå fast en europeisk vattenpolitik .
129 kemiska ämnen skulle regleras .
I slutändan fastställdes normer för endast ett tiotal ämnen .
Orsaken till det misslyckandet var enhällighetsprincipen .
För ungefär sju år sedan verkade det också som om den europeiska vattenpolitiken skulle offras på subsidiaritetsaltaret .
De konservativa regeringscheferna Major och Kohl beslutade vid toppmötet i Edinburgh att det inte alls var nödvändigt att spanjorer fick lika bra dricksvatten som tyskar och engelsmän .
Delvis tränger den inställningen igenom i den gemensamma ståndpunkt som tillkom under det brittiska socialdemokratiska ordförandeskapet .
Den ståndpunkten är en ost med hål i , eller för att använda vattentermer , den läcker som ett såll .
Det förklarar stormfloden av ändringsförslag från utskottet för miljö : nästan hundra ändringsförslag till den andra behandlingen .
Det är ovanligt att göra så men de flesta ändringsförslagen behövs verkligen för att täta alla läckor .
En stor läcka är de farliga kemiska ämnena .
Den kemiska industrin och tyvärr även Europeiska kommissionen och ministerrådet vill göra en enskild riskanalys för varje farligt ämne .
Det tar lång tid , och ännu viktigare , det finns ingen godtagbar nivå för föroreningar genom farliga kemiska ämnen .
Endast havets bakgrundsnivå är godtagbar .
Det är det som menas med termen " close to zero " .
Kommissionen har redan utarbetat en lista med 32 ämnen som prioriteras .
Många av dessa har en hormonstörande verkan .
Det är de så kallade endocrine disrupters .
De förorsakar till och med i ytterst minimala mängder könsförändringar hos djur och till och med hos människor , vilket ofta fastställts av vetenskapsmän .
Därför är det så viktigt att Europaparlamentet uttalar sig för Ospar-målet på nästan noll år 2020 .
Jag vill ta upp två av de ämnen som finns med på kommissionens lista .
Kvicksilver och tributyl , förkortat TBT .
På botten av Waddenzee ligger värdena för kvicksilver och TBT tio respektive tusen gånger högre än Ospar-värdet .
Den kemiska industrin och samhället som helhet måste lära sig att byta ut de här farliga ämnena mot oskadliga ersättningar , och om det inte går , att hantera dem i slutna system .
För medlet TBT betyder det att det inte längre får användas som medel för algbekämpning .
Mekanisk rengöring av fartygssidorna är ett bra alternativ .
Låt mig avsluta med att uttala min förhoppning om att Europaparlamentet hämtar upp sin gröna framtoning igen och uttalar sig för nästan noll-alternativet när det gäller farliga kemiska ämnen och hormonstörande ämnen till år 2020 .
Herr talman !
I behandlingen av detta direktiv om vatten har parlamentet en avgörande roll .
Rådets gemensamma ståndpunkt är helt otillräcklig inom flera områden .
Det måste därför nu vara vår uppgift att strama upp och konkretisera kraven i direktivet .
För oss i GUE / NGL-gruppen har några principer varit speciellt viktiga när vi har tagit ställning till de olika förslagen .
För det första anser vi att tidsramarna för att genomföra åtgärderna i förslaget måste bli kortare än vad rådet har föreslagit .
Vi stöder därför förslagen om snävare tidsramar för att genomföra olika delar av direktivet .
För det andra vill jag att utfasningen av farliga ämnen skall ske på ett konsekvent sätt .
Den får inte fördröjas av att man framför nya krav på utvärderingar innan åtgärder vidtas .
I lagstiftningen måste också respekten för internationella konventioner som Ospar-konventionen skrivas in .
För det tredje vill vi att prispolitiken skall vara klart uttryckt .
Det innebär att grundprincipen måste vara att man betalar de verkliga kostnaderna för vattnet .
I dag får skattebetalarna ofta subventionera industri och jordbruk .
Att förorenaren eller förbrukaren betalar skall vara den självklara utgångspunkten för lagstiftningen , även om det också kan krävas undantag i vissa extrema fall .
För det fjärde vill vi att undantagen från reglerna på vattenkvalitetområden skall vara få och tydligt avgränsade .
För det femte vill vi att skyddet av grundvattenkvaliteten och åtgärder mot fortsatta föroreningar i grundvattnet skall vara tydliga och klara .
Mot denna bakgrund kan vår grupp rösta för ett flertal av föredragande Lienemanns ändringsförslag , såsom de antogs i utskottet .
På ett par punkter skulle vi vilja gå ett steg längre .
Vi kommer därför att rösta för De grönas ändringsförslag 102 , 103 och 104 , som vi tycker ytterligare förbättrar positionen .
Vad gäller prispolitiken förekommer ibland extremsituationer , som kan kräva undantag från principerna i betänkandet .
Jag anser möjligheterna till undantag vara väl tillgodosedda i ändringsförslag 43 från utskottet och uttryckta på ett ännu bättre sätt i ändringsförslag 105 från De gröna .
Jag kan inte se att det skulle behövas några ytterligare undantag än de som anges i dessa två ändringsförslag .
Detta finns det emellertid olika meningar om inom vår partigrupp .
Ändringsförslag 107 , som berör frågan , har lämnats in av en del av vår grupp .
Som helhet tycker jag att förslagen från utskottet i Lienemanns betänkande är bra , och kan vara en god grund för en svår förlikning .
Herr talman !
Alla fotografier som tas av satelliter visar att vi verkligen bor på den blå planeten : detta vattenöverflöd är dock en illusion .
Den katastrof som nyligen inträffade i Donau påminner oss om att floder och älvar är jordens vitala artärer och att föroreningar inte har några gränser .
Vatten är en förnybar och begränsad naturresurs .
Det minskar då det inte förvaltas på rätt sätt och de geografiska och klimatiska förhållandena inte är gynnsamma .
Inom EU är detta en avgörande fråga i Medelhavsområdet , men också i andra länder i Europa , där vi ser en progressiv uttorkning av våtområden .
Känsliga , våta eller torra områden , olikheter mellan stater , olikheter mellan olika regioner inom staterna samt klimatiska , ekonomiska , geografiska , geologiska särdrag är i hög grad bevis som vi vill påminna om men som inte för den skull bör leda till snedvridningar av konkurrensen i gemenskapen .
Vi har dock ingett ändringsförslag för att påminna om betydelsen av jordbrukets specifika relation till vatten , en viktig faktor för markanvändning och -bearbetning .
Självklart är jordbrukets behov större i söder och detta särdrag måste beaktas i ramdirektivet .
Det är för övrigt inte bara i unionens stater som man söker lösningar på dessa problem : partnerskapsländerna i EU-Medelhavsområdet begärde i Turin i oktober en Marshallplan om vatten för Medelhavets södra kust .
Lyckligtvis är vi inte där ännu .
I Europa finns likväl torka , en ökenutbredning av vissa områden , men också översvämningar , och direktivet understryker detta .
Vi drabbades nyligen av det i Frankrike , också i Rhendalen och Centraleuropa .
Vi behöver detta ramdirektiv såsom en väsentlig beståndsdel av en hållbar utvecklingspolitik , som bör göra de olika användningarna av vatten kompatibla sinsemellan .
Men det är nödvändigt att man i denna nya förvaltning införlivar skydd och bevarande av den biologiska mångfalden .
Ärendet " vatten " kommer under alla förhållanden inte att avslutas i dag .
Frågan om utvidgningen och klimatförändringarna öppnar nämligen nya framtidsutsikter .
Herr talman !
Vatten av god kvalitet kommer det här seklet kanske att ha ett ännu större strategiskt värde än olja .
Det är skäl nog att tacka Lienemann för hennes insatser för att ytvattnet skall få en stark ställning .
Det verkar vara ganska invecklat att komma fram till en bra ram för den europeiska lagstiftningen .
Med ramdirektivet för vattenpolitik vill vi göra slut på den splittrade vattenlagstiftningen i unionen .
Därmed undkommer vi emellertid inte ett omfattande och komplicerat direktiv .
För det krävs att de verkställande instanserna är mycket noggranna vid genomförandet av det .
Särskilt viktigt är det att medlemsstater och vattenmyndigheter utnyttjar sina möjligheter att föra en specifik politik , som tillkommit tack vare tillvägagångssättet med avrinningsområden .
De viktigaste målen förblir att bekämpa en ytterligare nedsmutsning av grund- och ytvattnet , skydda ekosystemen , stimulera en hållbar användning av vatten , bekämpa översvämningar och torka samt att sluta släppa ut farliga ämnen i ytvattnet .
När det gäller utsläppen av farliga ämnen så anser jag att rådets målsättningar är för vaga och inte tillräckligt ambitiösa .
Förslaget från miljöutskottet att föra tillbaka utsläppen till nästan noll tycker jag är sympatiskt och eftersträvansvärt .
Det måste dock ägnas mycket uppmärksamhet åt genomförbarheten .
Därvid måste hänsyn tas till naturliga bakgrundsutsläpp som inte kan påverkas och även svårhanterliga diffusa utsläpp som ändå förorenar vattnet rejält .
Herr talman !
Vi måste under 2000-talet ta till oss den grundläggande tanken att vi har ett helt nytt förhållande till vattnet .
Under 1900-talet var vattnet för oss ett kostnadsfritt transport- och avfallssystem för gift , farligt avfall , kemikalier osv .
Följderna ser vi redan !
Vi måste tänka om och erkänna vattnet som vår viktigaste livspartner , och vårt ansvar för detta går långt utöver de nuvarande generationerna .
På så sätt måste också direktivet behandlas under förlikningen , och befolkningen måste kunna förstå vad vi här planerar , respektive vad kommissionen planerar .
Skyddet för vattnet är principiellt också en social fråga , och en avgörande sådan .
Därför skall principen " förorenaren betalar " användas i större utsträckning , eftersom följderna annars måste bäras av alla .
Med tanke på de långtgående skadorna på vattenresurserna är det viktigt att vi inte bara bibehåller nuvarande nivå , utan i morgon vid omröstningen ser till att det skapas verkliga kvalitetsförbättringar .
Herr talman !
Det är nu redan cirka sex år sedan som vår kollega Karl-Heinz Florenz , assisterad av Ursula Schleicher , bad om en omstrukturering av hela vattenpolitiken .
Det lyckades .
Det är inget enkelt ämne och jag tycker att de insatser som Lienemann gjort förtjänar stor respekt .
Beslutsfattandet kring det här ramdirektivet befinner sig i ett mycket viktigt skede .
Ämnet har förts in under medbeslutandeförfarandet och vid den första behandlingen har vi därigenom redan kunnat skapa en viktig och sträng lagstiftning .
Den gemensamma ståndpunkt som lades fram i slutet av förra året är också en viktig förbättring jämfört med det ursprungliga förslaget .
Det är också mycket svårt att föra en politik på den här punkten eftersom skillnaderna är så stora .
Till min spanska kollega säger jag : i norra Europa har vi ofta översvämningar att tampas med men även förorenat vatten från industrin , medan problemet för kollegerna i söder ofta är att vatten måste transporteras långa avstånd helt enkelt för att ge dricksvatten eller vatten för jordbruket .
Jag skall gå in på de två aspekterna av det här ämnet .
Först kvaliteten .
Nederländerna påverkas till stor del av den europeiska vattenpolitiken .
En mycket stor del , en tredjedel av vårt dricksvatten , utvinns i Nederländerna från ytvatten .
Nederländerna ligger nedströms , i ett delta , och därför är alltså kvaliteten på det ytvatten som kommer till oss av allra största vikt .
En annan viktig diskussionspunkt är normerna för vattenkvalitet .
I ett antal ändringsförslag sätts det frågetecken för de föreslagna normerna och särskilt med avseende på Ospar-normen för år 2020 .
Jag förstår väl att vissa tycker att den normen är otydlig eller juridiskt oförsvarlig .
Jag tycker dock att vi måste stödja den eftersom vi då kan ombesörja noggrannare normer i förlikningsförfarandet .
Sedan några ord om kvantitetshanteringen .
En berömd nederländsk poet talade redan i sin dikt " Minnen från Holland " om vattnet som fruktades på grund av de ständiga katastroferna .
År 1953 inträffade en jättelik vattenkatastrof , varigenom vi samtidigt även blev föregångare när det gäller fördämningar .
År 1990 svämmade våra floder över och vi kunde konstatera att anläggning av konstgjorda verk uppströms påverkar förmågan att ta emot vatten nedströms och kan leda till stora skador .
Det betyder att vi även när det gäller kvantitetshantering måste göra stora ansträngningar för att se till att det går bra att leva både uppströms och nedströms .
Herr talman !
Jag skulle gärna vilja börja med att ge Lienemann mina välmenta komplimanger .
Hon har gjort ett utmärkt arbete .
Vatten är ett första livsbehov och en grundläggande rättighet .
Var och en borde ha tillgång till rent vatten men tillgång och bra kvalitet på vatten är inte någon självklarhet , det får många erfara , i Sydeuropa men nu också i länderna längs Donau .
Vatten är ofta en källa till konflikter mellan länder och mellan befolkningsgrupper .
Därför är det viktigt att vatten blir föremål för internationell samordning .
Vi måste erkänna att vatten är vårt gemensamma ansvar .
Samarbete inom ett avrinningsområde måste vara en självklarhet .
För liten kapacitet uppströms eller just en för riklig användning kan skapa problem nedströms .
Samordning är nyckelordet här .
Vattenproblemet blir allt aktuellare .
Förändringar i klimatet , små temperaturhöjningar påverkar nederbörden direkt .
Vissa områden blir torrare , många områden blir våtare .
Det är dags att göra något .
I mars anordnas ett andra världsvattenforum i Haag .
Det här forumet står för en världsomspännande vision .
Den visionen måste leda till regionala handlingsplaner för hållbar förvaltning och hantering av vatten .
För Europaparlamentet har det nu blivit dags att handla .
Vi måste nu ta ställning för en hållbar vattenpolitik som utgångspunkt och samtidigt måste vi vara realistiska .
Vi får dock inte heller lägga ribban för lågt .
Den gemensamma ståndpunkten är inte tillräckligt ambitiös .
Därför är det nödvändigt att vi griper tag i tidigare internationella avtal eller Ospar-målen .
Vi måste sträva mot en utfasning av farliga ämnen år 2020 .
Det är redan avtalat för havsmiljön .
Det ligger nära till hands att det här avtalet även skall gälla för andra vatten .
Ospar-målen håller nu på att utarbetas .
Det har ställts upp en lista med 400 ämnen som innebär tydliga risker för miljön .
Både tekniskt och ekonomiskt är det genomförbart att i princip minska utsläppet av de här ämnena till noll och det måste vi nu ta ställning för igen .
Direktivet skall naturligtvis också vara bindande .
Länder nedströms måste kunna lita på att länderna uppströms uppfyller kvalitetsmålen .
Kvalitet har ett pris men förorening kan visa sig bli ett mycket högre pris att betala i framtiden .
Herr talman , fru kommissionär !
Jag vill uttrycka min djupa respekt för det utomordentliga arbete Lienemann utfört med detta vattendirektiv .
Låt mig påminna om att de riktigt stora miljöproblemen i dag - klimatförändring , skövling av urskogar , utfiskning av haven - hela tiden berör våra gemensamma och absolut nödvändiga , men på något sätt herrelösa resurser .
Låt oss också inse att vårt färskvatten i Europa kan sägas ligga i gränslandet mellan att ägas av alla och av ingen .
Därför är det strategiskt viktigt att ansvaret för vattnet fastställs .
Det är också viktigt att de olika vattendragen hålls samman och hanteras som den helhet som de är , oavsett vem som äger den ena eller andra delen av ett gemensamt vattenflöde .
Kära kolleger !
Förslaget till direktiv utgör i själva verket , som redan flera gånger sagts , en historisk möjlighet att förenkla och förbättra oredan och trasmattan av EU-förordningar och direktiv , och på så sätt uppnå en hög miljöskyddsnivå i Europa .
Men jag har fått det intrycket att vattenramdirektivets politik präglats av avreglering och åternationalisering .
Jag hoppas också att omröstningen inte blir till ett slag i vattnet , och därför är två punkter väsentliga för mig .
För det första Ospar .
Vi känner till att kommissionens förslag inte går tillräckligt långt ; tyvärr gäller detta också för förslaget från utskottet för miljö , folkhälsa och konsumentfrågor .
Att bara slumpmässigt lägga fram förslag , räcker inte .
Det vi behöver är ett rättsligt absolut bindande mål för Ospar .
Endast då kommer vi att kunna åstadkomma rättslig klarhet och framför allt möjligheter till överklaganden .
Allt annat skulle förfela sin verkan och inte bidra till att förhindra att ekologiska katastrofer , liknande dem som vi nu upplever i Rumänien och Ungern , också skulle kunna inträffa hos oss .
Jag finner det beklagligt att de nationella regeringarna inte är beredda att engagera sig för ett rättsligt bindande skydd , fastän de ju internationellt har enats om Ospar .
Men jag tror att det är just det som vi här i parlamentet måste ordna upp , för att därigenom visa att vi inte tillåter att vår trovärdighet utsätts för någon förlust eller någon skada .
Det som är viktigt är också att stärka principen om att " förorenaren betalar " , ty priserna måste säga den ekologiska sanningen .
Vi får inte ge efter för jordbruks- och kemiindustrins lobbyintressen , utan vi måste propagera och med vår omröstning ge uttryck för att vi vill ha principen " förorenaren betalar " och därmed få kostnadstäckande priser .
Vatten är den viktigaste resursen för vårt liv , och vi måste med vår omröstning se till att det finns impulser och påtryckningar för att verkligen iaktta Ospar-konventionen .
Med hjälp av slutna kretslopp i produktionen är detta möjligt , allt annat skulle vara en urvattning av direktivet .
Låt oss ta denna chans !
Herr talman !
På den korta tid jag har till mitt förfogande vill jag välkomna föredragandens betänkande och påminna om tre principer som bör vara överordnade de övriga , och som tydligt kommer till uttryck i föredragandens ändringsförslag : vattnet är inte en kommersiell produkt utan något som tillhör unionens folk ; det yttersta målet är att lyckas utplåna alla förorenande ämnen av ytvattnet och grundvattnet , och behovet av att informera befolkningen så att den kan medverka till att återvinna vattnet och inte slösa med det som är en så värdefull resurs .
Jag vet att det kan bli problem med det här direktivet , för man talar här om att verkligheten skiljer sig åt i unionens olika länder .
Det som händer i norr är inte det samma som det som händer i söder , inte heller som i de länder där man har problem med ökenutbredning .
Jag är medveten om det .
Men vissa ändringsförslag försöker hjälpa länderna i söder , närmare bestämt ändringsförslag 43 som , när det gäller att återvinna kostnaderna , även anger att medlemsstaterna bör ta hänsyn till ländernas sociala och miljömässiga villkor när beslut fattas .
Även överledningen av vatten är ett problem .
I mitt land - jag bor i norra Spanien - är det stora skillnader mellan norr och söder , och svårigheter uppstår när vattnet skall överledas från en plats till en annan .
Men det framgår även av Lienemanns betänkande att man i uppsamlingsplatserna bör spara på och värna om vattnet .
Jag är medveten om att det är ett komplicerat betänkande , att det finns olikheter beroende på de skilda verkligheterna i länderna , men vi bör föra fram ett ramdirektiv som förhindrar en upprepning av det som händer i Donau och det som hände i Doñana .
Vi kan inte tillåta att man förorenar Europas vatten , herr talman , och vi bör upprätta ett direktiv som förstärker regeringarnas politiska vilja att bevara en resurs som vattnet , som är så värdefull för alla .
Herr talman !
Jag gratulerar föredraganden till ett utmärkt betänkande .
Som irländsk ledamot av Europaparlamentet som kommer från ett land med stora vattenreserver stöder jag de stora flertalet av förslagen i detta direktiv .
Jag skulle emellertid nu vilka granska de sakfrågor som skiljer mellan parlamentets utskott för miljö och rådet .
Det senare har redan presenterat sin gemensamma ståndpunkt om denna fråga .
Enligt rådet skall målet att uppnå bra ytvattenstatus kunna uppnås senast 16 år efter det att direktivet träder i kraft medan parlamentets utskott för miljö vill få denna tidsfrist förkortad till tio år .
Jag ser inget skäl till varför Europeiska unionens medlemsstater inte är i stånd att genomföra de centrala bestämmelserna i detta direktiv under så kort tid som möjligt .
Jag övergår nu till de ändringsförslag som skall läggas fram för parlamentet i morgon om principen om omkostnadstäckning för vattenutnyttjande .
Rådet fastslår i sin gemensamma ståndpunkt att Europeiska unionens regeringar måste ta hänsyn till principen om omkostnadstäckning för vattenutnyttjande .
Inget bestämt slutdatum för att genomföra denna princip fastslogs i den gemensamma ståndpunkten .
Ändringsförslag 43 som innebär att man vill sträva efter att senast år 2010 kunna garantera att vattenprispolitiken i Europa skapar tillräckliga incitament för ett effektivt vattenutnyttjande .
Vidare skall ett adekvat bidrag från olika ekonomiska sektorer , uppdelat i industri- hushålls- och jordbrukssektorn , garantera att denna politik genomförs .
Om dessa ändringsförslag inte stöds i morgon kommer en stark signal sändas ut att mätare och vattenavgifter bör införas för hushåll i alla stater i Europeiska unionen .
Detta är politiskt opraktiskt ur irländskt perspektiv liksom det faktiskt skulle vara ur andra medlemsstaters perspektiv som Portugal , Grekland och Spanien .
Herr talman !
Först och främst vill jag gärna tacka Lienemann för hennes betänkande .
Det är här och nu vi avgör om EU-länderna skall arbeta effektivt för en renare vattenmiljö under de kommande åren .
Det gör vi som parlament genom att ändra rådets gemensamma ståndpunkt och visa den väg som leder fram till ett samarbete för en renare miljö .
I oförändrad form kan detta direktiv nämligen få mycket olyckliga och långvariga konsekvenser för miljön och dricksvattnet .
Det skulle innebära att man skickade fel signaler till både den europeiska industrin och den europeiska befolkningen .
Det är avgörande att stå fast vid en begränsning av det totala utsläppet av kemiska ämnen i våra vattenområden .
Det resulterar uppenbarligen i en alltför utdragen tidsaspekt om man skulle göra mätningar av varje enskilt ämne som finns i omlopp , eftersom det finns ca 100 000 .
Vi har inte råd att vänta .
I detta sammanhang ber jag parlamentet att stödja ändringsförslag 108 , där orden " förorening av vatten genom enskilda förorenande ämnen " , ersatts av " förebyggande av förorening av vatten genom att fortlöpande minska utsläpp " .
Vi kan inte försena miljöarbetet genom att överdriva detaljerna i stället för att verka för en minskning av de totala utsläppen av farliga ämnen i miljön .
Denna konvention skall vara en riktlinje i arbetet för den rena miljö som vi är skyldiga oss själva och inte minst våra efterkommande .
Herr talman !
Det är svårt att sammanfatta huvuddragen i ett direktiv som är så viktigt och komplicerat .
I Amsterdamfördraget slås fast att vi skall prioritera förebyggande åtgärder , tillämpa principen att " den som förorenar betalar " och skapa en hållbar utveckling där miljökonsekvenserna tas med i beräkningen .
Det är viktigt att man urskiljer det ekonomiska värdet av miljöpåverkan vid prissättning och får aktörerna att ta sitt ansvar genom att införa incitament att använda icke förorenande system .
Detta är odiskutabelt mot bakgrund av förhållandet mellan ekonomisk utveckling och tryggande av miljön , särskilt vattentillgången .
Denna situation tar sig specifika uttryck inom många ekonomiska sektorer , men särskilt inom jordbruket .
I det komplicerade förhållandet mellan jordbruk , miljö och vatten , mellan positiva och negativa konsekvenser , mellan en mängd olika lokala situationer och produktionssystem och så vidare , har man infört konceptet om god jordbrukspraxis .
Med detta avses den produktionsmetod som används inom jordbruket så att man uppfyller gemenskapens förväntningar på att man skall hålla vården av vattenresurserna på en högre nivå än minimistandarden , med därav följande kostnader och minskade intäkter .
Ur detta koncept härrör tvånget att bygga ut och förstärka en integrationsstrategi för att bibehålla vattenvården i centrum av den ekonomiska produktionsmodell som är hållbar mot bakgrund av gällande förutsättningar .
I ljuset av detta skall man inte följa strategin att skilja målsättningen att förhindra att yt- och grundvattnet försämras från målsättningen att skydda , förbättra och återställa dess kvalitet , och därmed skapa en konstgjord prioriteringsskala till förfång för en heltäckande insats med specifika riktade åtgärder inom ramen för denna och där man använder bästa tillgängliga teknik .
Vad beträffar att eliminera de föroreningar som härrör från farliga ämnen i vattenmiljön bör man för att optimera tillvägagångssättet införa bestämmelser på både nationell och gemenskapsnivå , så att man bättre kan identifiera de olika typer av vattendrag som förorenats till följd av människors produktion .
Slutligen måste man konstruera ett system som innehåller en objektiv förteckning över potentiellt farliga ämnen med mesta möjliga information om kemiska , fysiska och biologiska egenskaper , för att skapa en integrerad modell för insatser på olika strategiska nivåer till skydd för tillgången på vatten som är oundgänglig för oss alla .
Herr talman , fru kommissionär , kära kolleger !
Om vi tar principen om hållbarhet på allvar , vilken ju är fastslagen i Amsterdamfördraget , då kan vårt långsiktiga mål i själva verket bara bli att uppnå nollutsläpp i vårt vatten .
Ty vi måste naturligtvis säkra vattnet så att kommande generationer inte belastas av hur vi använder vattnet .
Därför gäller det här att utveckla steg med anspråksfulla normer , för att uppnå detta långsiktiga mål .
Därför stöder jag eftertryckligen Lienemanns ändringsförslag för att här utveckla en förnuftig väg med kvalitetsnormer , så att vi verkligen någon gång kan säga att mänsklig användning av vatten faktiskt inte betyder förbrukning av vatten , utan säkrar vattnet i det tillstånd det befinner sig .
Direktivet erbjuder några mycket positiva beståndsdelar , som absolut kan framhävas än en gång .
För det första är det den faktiskt breda informationen till allmänheten och delaktigheten för den .
Det har det knappast funnits i något europeiskt direktiv .
För det andra är det tvånget till samarbete .
Jag anser att det är glädjande att man här betraktar vattenresurserna som en helhet och att myndigheter , både i de enskilda medlemsstaterna men också utanför medlemsstaternas gränser , äntligen tvingas samarbeta och se till att det blir en hög nivå på kvaliteten i samtliga vattenresurser .
För det tredje vill jag också ta upp frågan med tidtabellen .
Jag är fullständigt övertygad om att vi behöver en strikt tidtabell , så att det också görs ansträngningar för att vi skall nå vårt långsiktiga mål .
Jag vill gärna jämföra det med situationen i december .
I december vet vi alla att det är jul den 24 , och vi börjar köpa julklappar .
Men hur vore det om vi i december visste att julen skulle inträffa om trettio år ?
Vi vet alla hur vi då skulle bete oss .
Därför behöver vi just när det gäller vattenpolitiken en strikt tidtabell .
Jag stöder eftertryckligen föredragandens förslag och anser att vi för alla områden i detta direktiv - vare sig det är en åtgärdslista eller frågan om sysselsättningsåtgärder - behöver en strikt tidtabell .
Herr talman !
Syftet med detta direktiv bör vara att se till att medlemsstaterna genomför samlade åtgärder för skydd av grund- , dricks- och ytvattnet , och att skyddsnivån motsvarar bestämmelserna i den befintliga gemenskapslagstiftningen på miljöområdet .
Låt mig här påminna om att tidigare beslut om nitratdirektivet ännu inte genomförts i samtliga medlemsstater , trots att det är ett gemensamt EU-beslut .
Detta förslag innehåller en rad åtstramningar av skyddet för vattenmiljön , som går utöver vårt nuvarande miljömål .
Det föreslås att man skall uppfylla ett slutmål för koncentrationer i havsmiljön nära bakgrundsvärdena för naturligt förekommande ämnen och nära noll för syntetiska ämnen skapade av människan .
Det är omöjligt och dessutom naturvidrigt .
Antagandet av detta betänkande kommer att få allvarliga konsekvenser för jordbruksnäringen i EU , om koncentrationen av t.ex. fosfor och kväve inte får överstiga bakgrundsvärdena för dessa ämnen i vattenmiljön och om man kommer att fastställa ett nollgränsvärde för bekämpningsmedel i vattenmiljön .
Jordbruket i Europa kommer t.ex. inte att kunna odla brödsäd med förhöjt proteininnehåll , så att säden kan användas till bröd .
Resultatet kommer att bli att jordbruksproduktionen flyttar till andra länder utanför EU , med stora sysselsättnings- och samhällsekonomiska kostnader som följd .
Jag kan inte rösta för de avsnitt i vattenramdirektivet som behandlar dessa förhållanden .
Herr talman , ärade kolleger !
Vatten är en dyrbar råvara .
Miljoner människor har inte ens tillgång till rent vatten , ett absolut villkor för att överleva .
Vi behöver därför inte förundra oss över att vatten ofta är en orsak till krig .
Den kapitalistiska världen placerar också ut sina spelpjäser för att få maximal kontroll över vattenförråden .
Därvid är det sällan tal om något allmänintresse eller någon solidaritet .
Europa står alltså inför en svår uppgift : föra samman den , både när det gäller mål och medel , splittrade vattenpolitiken i gemenskapen i en mer sammanhängande ramlagstiftning .
Jag måste bekänna att även i mitt land , Flandern , är det en lång väg att gå .
Även vi fick nyligen smäll på fingrarna av kommissionen för det .
Varje förnuftig människa vill att det här ramdirektivet används som ett påtryckningsmedel för de politiska ledare som nu kommer till korta .
Den gemensamma ståndpunkten är i det avseendet en fars , ett verk utan tvång , en riktig förolämpning mot Ospar-avtalen .
Vi har till och med en tidsfrist för genomförande som kan tänjas ut till 34 år framåt .
Mina barn kommer då att vara äldre än vad jag är nu .
Håll med om att det här inte är rätt .
I morgon kan vi välja en svag ram utan tvångsmekanism som förgiftar framtiden för våra barn .
Antingen röstar vi för ändringsförslagen från min grupp , från föredraganden eller från utskottet för miljö .
Bara en sak till .
De senaste månaderna har det varit en enorm lobbyverksamhet på gång .
Vad som var iögonenfallande i den här saken var den enorma pressen från ministerrådet .
I mitt eget land skedde det både genom de flamländska och de wallonska miljömyndigheterna .
De ställer sig bakom den svaga gemensamma ståndpunkten till förmån för ett ytterligare ställningstagande av vårt parlament .
Jag undrar verkligen om det här är ett försök som de gröna miljöministrarna i mitt land känner till .
Kolleger !
Det räcker inte längre med vackra ord .
Vi måste göra en resolut kursändring .
Vid omröstningen i morgon kan vi göra det tydligt att Europa anstränger sig för att skapa en ansvarsfull och framtidsinriktad vattenpolitik .
Det kan bara öka vår trovärdighet .
Jag förklarar debatten avbruten och den kommer att återupptas kl .
09.00 .
 
Dialog om Europa : institutionella reformens insatser Nästa punkt på dagordningen är kommissionens meddelande - Dialog om Europa - institutionella reformens insatser .
Herr talman , mina damer och herrar ledamöter !
I kommissionen pågår just nu en debatt och mycket skall till för att detta arbete skall avslutas i dag .
Jag kommer huvudsakligen för att , såsom angetts på föredragningslistan , tala om ett nytt initiativ som kommissionen förslår till svar , och det är inte det enda svaret , på en stor utmaning som bör mobilisera samtliga aktörer i den europeiska uppbyggnaden , i vilken ni befinner er i första ledet i egenskap av parlamentsledamöter , men också jag såsom kommissionsledamot , också de ministrar som sitter i rådet , de nationella parlamentsledamöterna och jag vill tillägga till och med de tjänstemän som arbetar i de olika institutionerna och som är engagerade i och motiverade av denna europeiska uppbyggnad .
I den långa debatten i morse där jag deltog vid sidan om ordförande Prodi berörde många av er det demokratiska underskottet och det stora avståndet till de europeiska institutionerna .
När jag säger det försöker jag inte bara att ställa frågan - en av er sade det mycket tydligt och med stor kraft : vem gör vad ?
Och det minsta man kan begära är att medborgarna förstår vem som gör vad i våra olika institutioner .
Frågan ställs då omedelbart också om vad vi gör tillsammans och vad vill vi göra tillsammans i framtiden , i synnerhet med de länder som skall ansluta sig till oss .
Det demokratiska underskottet får oss således också att undra och därför beslutade vi nyss i kommissionen att redan dagen efter öppnandet av regeringskonferensen , under vilken jag har fått äran att företräda kommissionen vid Prodis sida , och i nära samarbete med era båda företrädare , Brok och Tsatsos , lägga fram " En dialog för Europa och om Europa " och att för vår del delta i direktkontakten med medborgarna .
Samtliga kommissionsledamöter har åtagit sig att varje gång som de måste bege sig till ett land , och inte bara sitt ursprungsland , och till ett område - för min del händer det tre eller fyra gånger per månad - ägna ett ögonblick av sin tid åt en direktdialog med medborgarna , inte bara med eliten eller de institutionsansvariga som man vanligen möter utan också skapa en direktkontakt i ett universitet , ett gymnasium eller en fabrik , att söka kontakt med människor , svara på frågor och lyssna .
Det kommer att bli den del som vi tar på oss , såsom ni kommer att göra det själva när det gäller denna nödvändiga ansträngning och angelägna förpliktelse som består i att minska det demokratiska underskottet , det vill säga avståndet till medborgarna i förhållande till vad vi gör .
Vi vill att detta initiativ skall skötas i samarbete med medlemsstaterna och i förbindelse med Europaparlamentet .
Vi kommer att göra en regelbunden sammanfattning så att den allmänna opinionen mäts och man kan justera eller omorientera .
Vi vill också agera i samråd med de nationella parlamenten , de lokalt folkvalda , icke-statliga organisationer , arbetsmarknadens parter och media .
Opinionsnätverk , politiska grupper och partier , Europaparlamentets ledamöter , nationella parlamentsledamöter , folkvalda , det sade jag just lokala myndigheter eller nationella parlament , Regionkommittén , Ekonomiska och sociala kommittén , det civila samhällets organisationer och universitetsmiljöerna kommer att beröras .
Jag vill för övrigt påminna om - behöver jag göra det - att Europaparlamentet själv redan tog initiativet den 1 februari , och jag vill åter tacka ordförande Napolitano för det , att ordna ett första arbetssammanträde med företrädarna för de nationella parlamenten , det vill säga företrädare för medborgarna i varje stat .
Kommissionen kommer att föreslå medlemsstaterna att ansluta sig till denna åtgärd , antingen inom ramen för ett tillfälligt samarbete eller i ett mer strukturerat partnerskap .
Vi upprättar en plan för media och nära kontakter med EU : s ordförande och Europaparlamentets talman .
Jag har sagt på vilket sätt kommissionsledamöterna kommer att delta vid möten och besök ute bland människor .
Vi vill ha medborgardebatter .
Kan jag bara , utan att föreläsa - framför allt inte - och inte heller ge råd , påminna om att när jag hade äran att vara minister för Europafrågor i mitt eget land , kände jag behovet av att få en direktdialog med medborgarna och när jag varje vecka förde den dialogen direkt i olika områden upptäckte jag att det fanns ett enormt behov av att ge ett ansikte åt Europeiska unionen och jag åkte således med en ledamot från Europeiska kommissionen , inte bara de franska kommissionsledamöterna för övrigt , ambassadörer i tjänst i Paris , ledamöter från Europaparlamentet , och förde en dialog och jag upptäckte att det fanns oändliga frågor , att de var intelligenta , att människorna hade ett behov av att respekteras , att man lyssnade till dem och förklarade för dem .
Det är vad vi skall göra med stöd av ett budgetanslag på omkring fyra miljoner euro som vi ber er ställa till vårt förfogande .
Det kommer att bli nödvändigt att förhandla fram ett anslag inom ramen för budgeten år 2001 för vi vill föra fram och leda denna idé inte bara försöksmässigt , utan varaktigt år 2000 och 2001 , det vill säga under hela förhandlingen i regeringskonferensen och ratificeringsprocessen .
Vi kommer att inleda denna dialog i Bryssel den 8 mars i närvaro av sjuhundra unga provanställda i kommissionen .
Er talman , Nicole Fontaine , har accepterat att stå vid ordförande Prodis och flera kommissionsledamöters sida för att inleda den första dialogen och , mina damer och herrar ledamöter , jag kommer att se till att varje gång en kommissionsledamot inleder en dialog skall de ledamöter från Europaparlamentet som finns närmast tillgängliga kunna vara närvarande själva och ge sin synpunkt och förklara Europaparlamentets arbete och roll .
Ja , det var vad jag ville säga , herr talman .
Jag är för övrigt beredd att svara på frågor , ta emot idéer och förslag från de ledamöter som är här .
Kolleger , ni känner till bestämmelserna .
Ni förväntas ställa frågor och inte nödvändigtvis göra långa uttalanden .
Ni har en minut var att ställa er fråga .
Herr talman !
Jag vill ge uttryck för min och , tror jag mig kunna säga , utskottets för konstitutionella frågor , vars ordförande jag är , uppskattning av detta initiativ från kommissionen .
Detta initiativ motsvarar för övrigt de anvisningar parlamentet självt gav i sin resolution från den 18 november .
Jag har också hört de preciseringar kommissionär Barnier gav om förhållandet med och kopplingen till Europaparlamentet när detta program utformades .
Om ni tillåter kommissionär Barnier , skulle man inte i meddelandetexten kunna säga någonting mer om detta än den enkla , litet kalla , frasen " elle sera conduite en liaison avec le Parlement européen " ?
Jag tycker att det vore bra om man kunde betona denna överensstämmelse i avsikter och bemödanden , även eftersom jag kan urskilja ett speciellt samordningsproblem som är just det mellan kommissionens initiativ , som verkligen inte bara riktar sig till ledamöter i Europaparlamentet utan även till ledamöter i nationella parlament och vårt utskotts program .
Efter den studiedag den 1 februari som kommissionär Barnier hänvisade till och där kommissionens betydande bidrag var till stor nytta är vår avsikt att ta upp regeringskonferensens utveckling vid alla våra möten .
Vi kommer därför att ha ledamöter i de nationella parlamenten närvarande vid alla våra möten , ett kvalificerat och bestående deltagande hoppas vi , och detta kommer att bli en kanal som blir ett bra komplement till dem i kommissionens initiativ .
Tack , ordförande Napolitano , jag bekräftar att det vi föreslår överensstämmer fullt ut med andan i resolutionen av den 18 november och jag vill också här säga att jag har kunnat föreslå kommissionen detta initiativ tack vare min kollega Vivianne Redings samarbete och goda samförstånd samt att det genomförs i förbindelse med Günther Verheugen , eftersom allt som står på spel och de stora utmaningarna , som vi måste förklara och våra landsmän i varje land undrar över och frågar om , gäller både utvidgningen - utvidgningens möjligheter och risker - och den institutionella reformen .
Jag har mycket väl förstått er oro , ordförande Napolitano , och det kommer att bildas en interinstitutionell arbetsgrupp ( det första sammanträdet kommer att äga rum i mars ) .
Jag skall se till att vi går bortom det som litet torrt står i kommissionens text , att vi talar om mer än förbindelse , om gemensamt arbete och att man sålunda under dessa två år kan samordna de initiativ som ni tar och som vi tar , var och en å sin sida , men som vi tar tillsammans .
Mina damer och herrar ledamöter , låt mig säga att om vi vill inleda denna dialog finns det arbete för alla .
Herr talman , herr kommissionär !
Det är ljuv musik för mina öron att höra er nämna ordet medborgare så ofta .
I detta parlament talar man mer och mer om den allmänna opinionen : rädsla för allmänna opinionen , det är som ni vet litet paternalistiskt , men vårt parlament är nu en gång så och vi måste acceptera det .
Jag ville ställa en exakt fråga till er inom ramen för frågan om regeringskonferensen : jag tror mig veta att domstolen i Luxemburg håller på att noggrant behandla en viktig fråga som handlar om bedrägeribekämpning och OLAF .
Såsom ni vet finns det förvisso problem som berör parlamentet men också europeiska tjänstemän , för de är också europeiska medborgare .
Jag ville fråga er med tanke på hur brådskande denna fråga har blivit om kommissionen har tänkt på möjligheten att ändra struktureringen av organisationen för bedrägeribekämpning fullt ut genom att tänka ut en lösning som innebär att bedrägeribekämpning i medlemsstaterna liksom i de europeiska institutionerna skulle ingå i domstolens behörighetsområde .
Herr Dupuis , först och främst sätter jag stort värde på ordet medborgare i mitt offentliga liv .
Det är ett av de finaste orden i en demokrati och jag tror att det måste användas .
Vi skall föra en dialog med medborgarna , inbegripet med de anspråkslösaste eller med de människor som är längst bort ifrån besluts- och informationscentrerna .
Eftersom ni talar om regeringskonferensen vill jag bara med anledning av frågan om bedrägeribekämpning i synnerhet - om det nu handlar om att kämpa mot bedrägeri mot gemenskapens intressen och budget - påminna om att vi för övrigt i kammarens arbetsanda och kanske genom att gå samma väg , kan jag säga att vi tagit fasta på idén i kommissionens förslag om att inrätta en speciell och ny tjänst såsom europeisk åklagare ; denne skulle således ha befogenhet enligt fördraget , således av medlemsstaterna , att från början till slut undersöka ett ärende som eventuellt ifrågasätter gemenskapens intressen och budget .
Vi noterar helt klart och nästan kliniskt att det rättsliga samarbetet inte längre räcker till , inte räcker för närvarande för att effektivt kunna bekämpa dessa bedrägerier , var de än kommer ifrån , inifrån eller utifrån , och därför har vi lagt fram detta förslag om att inrätta tjänsten som europeisk åklagare , som efter att själv ha undersökt ett ärende från början till slut skulle kunna låta det undersökas därefter och dömas av lämpligaste nationella domstol .
Vi har inte - jag svarar på den andra punkten om domstolen - vi har ännu inte klargjort våra ståndpunkter om domstolen eftersom vi väntade på betänkandet Dur som inlämnades för några dagar sedan .
Såsom jag hade åtagit mig skall kommissionen komplettera sina förslag rörande yttrandet om regeringskonferensen , i fråga om domstolssystemet och domstolen , inom de närmaste veckorna .
Herr talman , herr kommissionär !
I förrgår visades en toppnyhet i det mest sedda danska nyhetsprogrammet , som jag vill be er kommentera .
Historien handlade om att en tjänsteman i kommissionen skulle ha sagt till en företrädare för det österrikiska näringslivet att eftersom han var österrikare så kanske han skulle utestängas från deltagande i ett vetenskapligt utbytesprojekt tillsammans med företag i andra länder , inklusive Danmark .
Jag vill be er att bekräfta att om en tjänsteman har sagt att ett österrikiskt företag på något sätt skall utestängas från deltagande i gemensamma utbytesprojekt , så har denna tjänsteman uttalat sig på ett felaktigt sätt , och om han inte har sagt så finns det ingen historia .
Kan ni bekräfta det ?
Herr Haarder !
Enligt min vetskap har ingen tjänsteman fått tillstånd att säga något liknande .
Det skulle inte vara , här uttrycker jag min personliga åsikt , normalt och rättvist att straffa de österrikiska medborgarna , företagen och de anställda på grund av oro över att en ny koalitionsregering bildats i detta land .
Med reservation för en kontroll som jag skall göra eller låta göra omedelbart efter sammanträdet bekräftar jag således vad jag sade : kommissionen har aldrig sagt eller beviljat något i den stilen .
Herr Haarder , det finns annat som vi rent allmänt kan lära oss av det som händer i Österrike .
Jag har själv tagit upp olika möjliga svar på denna utmaning som för oss alla består i att påminna om och att på nytt visa vad vi gör tillsammans sedan 1957 : en ekonomisk gemenskap , naturligtvis , men först och främst en värdegemenskap och en stadga om grundläggande rättigheter som kommer att mer och tydligare skydda enskilda medborgare , artikel 13 i fördraget rörande diskrimineringar .
Vi föreslog redan före den österrikiska krisen i vårt yttrande av den 26 januari att denna artikel efter regeringskonferensen skall omfattas av kvalificerad majoritet och inte längre av enhällighet , och det finns en eventuell möjlighet , jag säger eventuell , - det säger jag personligen - att komplettera artikel 7 med en ny strecksats som skulle förse förfarandet med övervakning eller demokratiskt larm på rättslig grund och sedan slutligen offentlig debatt .
Det enda sättet att få bort dåliga idéer är att ersätta dem med nya .
Jag återvänder därmed till ämnet för diskussionen : just nu tror jag djupt på debattens demokratiska värde och kraft , i synnerhet för att bekämpa demagogi .
Kommissionär Barnier !
Ni lade stor vikt i er redogörelse vid hur viktigt det är med en dialog med Europas medborgare .
Med hänvisning till regeringskonferensen , som ni vet , tilldelades enligt besluten i Helsingfors det portugisiska ordförandeskapet en speciell rätt att utöka dagordningen för konferensen under konferensens gång .
Utan tvivel har parlamentet sina egna företrädare , Brok och Tsatsos , närvarande .
Men kan ni , herr kommissionär , även lämna ett löfte att om och när dagordningen utökas av rådet så skall ni meddela detta till parlamentet så att vi kan diskutera det mellan oss själva och naturligtvis med er med avsikten att fortsätta den dialogen med medborgarna som ni lagt så stor vikt vid ? .
( FR ) Herr Beazley !
Mitt svar är ett klart och tydligt ja , men det är uppriktigt sagt ingen nyhet .
Ordförande Napolitano , många ledamöter från utskottet för konstitutionella frågor och ännu fler ledamöter här i plenarsammanträdet vet att jag kommer att vara tillgänglig för att under hela förhandlingen på kommissionens vägnar tala om hur det går i en anda av öppenhet och på realtid .
Jag kommer kanske att säga det på annat sätt än professor Tsatsos och Elmar Brok som är era direkta företrädare .
Det är för övrigt troligt att vi kommer att säga det tillsammans vid många tillfällen .
Jag tror att det är viktigt att förhandlingen inte är hemlig vare sig för Europaparlamentet eller för de nationella parlamenten , vilka , vill jag påminna om , i sista hand måste avge sin åsikt och inta en ståndpunkt i ratificeringsprocessen .
Därför hyllade jag Napolitanos initiativ till ett gemensamt och regelbundet samråd mellan de femton ländernas nationella parlament och Europaparlamentet .
Därmed börjar öppenhets- och debattskyldigheten här när det gäller institutionsreformen .
Jag kommer således att vara tillgänglig varje gång ni önskar det för att redogöra för våra ståndpunkter och framstegen i förhandlingen under hela detta år .
Herr talman !
I första hand mina komplimanger för kommissionens handlingssätt .
Jag tror att det är mycket bra att man inleder samtal med medborgarna i ett tidigt skede , det skedde ju inte vid Amsterdamfördraget eller vid Maastrichtfördraget och det har bara lett till en stor misstro .
Två frågor : för det första , ni har sagt att ni skall samtala med medborgarna och jag börjar redan med 700 praktikanter vid Europeiska kommissionen .
Tänker ni också rikta er till medborgarna via media , alltså även via TV och via Internet ?
Min andra fråga är en kritisk fråga .
Det har nyss lagts fram ett förslag om öppenhet och insyn från Europeiska kommissionen .
Om jag jämför det med det förslag som gäller för lagstiftning hos oss i Nederländerna så är det bara en liten skugga av det och det förslaget har lett till mycket kritik i Nederländerna .
Min fråga är egentligen : hur vill ni utforma öppenheten med avseende på regeringskonferensen , det direktiv som nu lagts fram är nämligen inte något bra exempel på det .
Fru ledamot , fru minister Maij-Weggen , eftersom vi talar om öppenhet när det gäller regeringskonferensen vet ni hur det kommer att gå till .
Förhandlingen börjar för övrigt just i detta ögonblick .
Representantgrupperna har sammanträde i Bryssel och jag skall skynda mig till dem strax .
Dokumenten kommer för det mesta att vara öppna , arbetsdokument .
Vi kommer inte att diskutera inför media under förhandlingssammanträdena som kommer att pågå under hela året mellan ministrarna och Europeiska rådet men jag har åtagit mig , jag kan inte göra annat just nu , att genomföra denna öppenhet och att redovisa i institutionerna om förhandlingen och om kommissionens ståndpunkt .
Jag vill bekräfta , samtidigt som jag tackar er för att ni frågat mig om det , att vi kommer att använda alla moderna medel , i synnerhet television , för att sända de offentliga debatterna i det ena eller andra landet , och till och med på europeisk nivå .
Vi kommer att öppna ett forum på Internet och skapa permanenta fora för diskussioner .
Kommissionsledamöterna skall åta sig att snabbt svara på alla frågor som ställs .
Vi kommer att använda alla dessa moderna medel .
Men jag tror att vi också måste anstränga oss att gå så nära inpå människorna som möjligt .
Jag skulle vilja att i samtliga Europas regioner - det är utan tvivel ännu litet utopiskt - skall en kommissionsledamot , när han kan det , en ledamot från Europaparlamentet , eller en minister kunna gå till offentliga debatter .
Jag har bevis för att det är möjligt .
De flesta av er gör dessa debatter i era valområden och i era regioner .
Ur kommissionens mer egoistiska synpunkt skulle jag vilja att denna institution får ett ansikte i medborgarnas sinnen och att de män och kvinnor som utgör den skall så ofta som möjligt kunna gå medborgarna till mötes .
Herr talman !
Jag uppskattar Barniers löfte att gå ut till regionerna , både för att förklara och för att lyssna till vad medborgarna har att säga .
Jag skulle vilja inbjuda honom till min egen region , Yorkshire , en större europeisk region som är en fullvärdig deltagare på den europeiska inre marknaden och en mycket stor mottagare av europeiska strukturfonder .
Han kan komma med båda de hattar han bär som en kommissionär .
Jag skulle vilja fråga honom hur energiskt kommissionen kommer att satsa på denna informationskampanj ?
I några medlemsstater är det inte bara fråga om att tillhandahålla information till en allmänhet som inte är så välinformerad som den kunde vara .
Det är naturligtvis viktigt men det gäller också att bekämpa den felaktiga information som sprids av en mycket aktiv anti-europeisk rörelse och av de anti-europeiska organisationer som finns .
Kommissionen måste ge mycket kraftfulla svar på några av de synpunkter som den kommer att få ta emot som en del av kampanjen .
Herr Corbett , jag tackar er för er uppskattning .
Jag accepterar gärna er inbjudan och om jag har förstått rätt , vill ni att jag , när jag kommer till Yorkshire , inte bara tar upp reformen av de europeiska institutionerna utan också strukturfonderna .
Jag kommer således att besöka er för att genomföra denna dubbla uppgift .
Jag glömde för övrigt att tala om hur angelägen jag är att möta , och jag har redan gjort det , de nationella parlamenten , inte bara genom att träffa deras företrädare här , utan genom att åka och träffa dem på plats .
För tio dagar sedan var jag i Westminster .
Ni ser , herr Corbett , att jag inte är rädd för svårigheter .
Jag skall nästa vecka besöka Bundestag i Berlin .
Jag har varit inför den franska senaten .
Under hela denna debatt kommer jag således att också varje gång det är möjligt direkt besöka de nationella parlamenten .
Vad beträffar dialogen med medborgarna handlar det inte om att göra propaganda eller marknadsföring , inte ens kommunikation .
Jag skulle vilja att dialogen verkligen blir en dialog , och att efter en liten film som objektivt förklarar vad som står på spel i fråga om den institutionella reformen , skall de som är här på tribunen kunna uttala sig och svara direkt .
Vi skall , jag upprepar det , genomföra detta initiativ till dialog i tillfälligt eller strukturerat samarbete med medlemsstaterna och jag vill mycket gärna med ert stöd att de femton medlemsstaternas regeringar skall kunna ansluta sig på de sätt som de anser lämpliga och passande till detta initiativ till dialog .
Herr talman !
Jag vill gärna ansluta mig till Barniers diskussionsgrupp med de 700 provkandidaterna , så han har några att diskutera med .
Det är ju inte så roligt att bara diskutera regeringskonferens och öppenhet med sig själv .
Under framställningen i parlamentet sade Barnier , i samband med regeringskonferensen , att socialpolitiken inte var underställd majoritetsbeslut , men när jag tittar på sidan 63 ser jag att kampen mot olika behandling , rätten att resa och att bosätta sig - alltså bosättningsdirektiven - hela socialförsäkringen , förnyelsen av förordning 1408 , av åtgärder på det socialpolitiska området - med ett fåtal undantag - skall underställas majoritetsbeslut .
Förstår inte Barnier att han går inte i hjärtat av medlemsstaternas valförfaranden ?
Det är ju p.g.a. dessa frågor som folk går till val och som leder fram till en ny majoritet i folketing och andra parlament .
Kan det styras från Bryssel ?
Är det ett led i den genomgripande decentralisering som Prodi talade om i förmiddags ?
Jag blev mycket glad när jag hörde förra veckan att kommissionen under flera år noga skall granska begreppet subsidiaritet avseende inte bara förbindelserna mellan union och medlemsstater utan också union , medlemsstater , regioner och städer .
Jag hoppas att kommissionär Barnier i sin strävan efter dialog i Europas regioner kommer att utveckla den tanken och lära av det han får höra .
Herr kommissionär !
Jag hänvisar till ett av era svar på de föregående frågorna där ni nämner det som jag kallar låsningen av fördraget inför snedvridningsriskerna , i synnerhet den mångfalden av sanktioner som kan drabba en medlemsstat genom tillämpning av artikel 7 för brott mot grundläggande fri- och rättigheter .
Tror ni att dessa förslag , eller förslag av denna typ , kan ingå i regeringskonferensens uppgift såsom den definierades i Helsingfors ?
Jag har för min del inte det intrycket .
Är ni inte rädd för att sådana sanktioner skall kunna slå slint och användas till att straffa , inte brott mot mänskliga rättigheter , utan små skiljaktigheter , åsiktsförbrytelser eller åsiktsskillnader i förhållande till den dominerande europeiska tanken ?
Ja , herr Bonde , vi kommer att inleda debatten med sjuhundra ungdomar i Bryssel .
Det är så att de kommer att arbeta i institutionerna och hos kommissionen och jag tror att det är bra att inleda debatten med ungdomar som är motiverade .
När det gäller det sociala trygghetssystemet vill jag bekräfta att vi har lagt fram förslag på området för kvalificerad majoritet eller på området för enhällighet utan ideologi .
I ert land , Bonde , liksom överallt tror jag att man är angelägen om att den inre marknaden skall fungera bra på de mest rättvisa villkor för konkurrens och rörlighet för varor och personer .
Och det är således det som är vår regel .
Vi föreslår nämligen att vi skall besluta med kvalificerad majoritet om vissa politiska områden , vissa skatteåtgärder eller i fråga om social trygghet och hälsovård när det har ett direkt samband med den inre marknadens funktion .
Vårt förslag är inte övergripande och det är inte systematiskt .
Jag känner mycket väl till hur känsliga dessa frågor är om beskattning och social trygghet .
Jag tror inte att vi skall stöpa samtliga nationella system för social trygghet i samma form , det har aldrig varit fråga om det , utan helt enkelt att säkra bästa villkor för den inre marknadens funktion i ett Europa med trettio eller tjugosju länder utan att en stat skall kunna låsa de tjugosex eller tjugosju övriga staterna .
Herr MacCormick , ja , jag bekräftar att denna dialog bör gå utanför de nationella huvudstäderna och att den bör gå så nära inpå människorna som möjligt , där de bor och har sina rötter och om jag sade något annat skulle jag inte vara överens med mig själv i egenskap av kommissionär med ansvar för regionalpolitik , det vill säga ett av de konkretaste och synligaste politikområdena , som är gjort för att stödja sysselsättning och livskvalitet för människor i regionen och ni kommer ofta att få höra mig säga att denna politik inte bara har skapats för det prioriterade målet med sammanhållning och solidaritet mellan regionerna , den har också skapats såsom ett komplement för att människorna skall kunna behålla sina rötter , sina traditioner , sin själ och sin identitet där de bor .
Vi skall således föra denna dialog med städer och regioner .
Berthu , Helsingforsmandatet är klart och tydligt och vi är inom denna ram .
Där planeras att de tre grundläggande ämnena som åsidosattes i Amsterdam skall behandlas först och prioriteras .
Tillhörande institutionella frågor läggs till samt slutligen frågor som det kan bli lämpligt , beroende på de portugisiska och franska ordförandeskapen , att tillföra under förhandlingen .
Kommissionen spelar sin roll om den tror att den bör komplettera i den ena eller andra frågan sitt yttrande som behandlar många institutionella frågor .
Jag är ännu inte säker på att vi kommer att göra det om artikel 7 och om vi gör det kommer vi inte bara att göra det till svar eller reaktion på en konjunktursituation , som är tillräckligt allvarlig för att de fjorton regeringarna i unionen har mobiliserats tillsammans för att lämna sitt svar och vi kommer också att göra det med tanke på framtiden i allmänhet .
Alla medel som definitivt kan stärka den värdegemenskap som vi utgör tillsammans alltsedan unionen grundades 1957 och till och med tidigare på ruinerna av andra världskriget , allt som kan göras kommer att vara lämpligt .
Herr Berthu , jag är säker på att vi kommer att kunna bli överens , ni och jag , på denna grund .
Tack , herr kommissionär .
Ni har besvarat frågorna noga och även inlett den dialog om Europa som hänvisade till .
Ni har visat ett mycket gott exempel på hur man håller tiden i dag .
Det avslutar debatten .
 
Frågestund ( kommissionen ) Nästa punkt på föredragningslistan är frågor till kommissionen ( B5-0009 / 2000 ) .
Första delen Fråga nr 36 från ( H-0025 / 00 ) : Angående : Hög barnadödlighet i Kosovo Enligt Världshälsoorganisationens senaste uppgifter till FN har Kosovo högst barnadödlighet i Europa ; nästan 50 procent av alla för tidigt födda barn dör .
Till följd av kriget har missfallen ökat kraftigt och de barn som inte föds för tidigt är mindre utvecklade än normalt .
Kan kommissionen , mot bakgrund av den humanitära hjälp som EU tillhandahåller och det politiska sändebudet Bernard Koushners ansträngningar , meddela vilka åtgärder den har vidtagit till skydd för kvinnorna i Kosovos rätt till moderskap och för gravida och födande kvinnors samt spädbarns hälsa ?
Herr talman !
Kommissionen är medveten om den mycket svåra situationen i fråga om hälsovård och hälsovårdsanordningar i Kosovo , inte bara för gravida kvinnor utan på hela fältet .
Detta beror både på den senaste konflikten och på alla år före konflikten av misskötsel och brist på underhåll .
Den statistik som nämns i fråga om barndödlighet talar för sig och är helt oacceptabel .
Situationen är dock knappast bättre för andra delar av befolkningen .
Kommissionens svar har varit följande : först och främst har hälsosektorn fått motta betydande bidrag från ECHO .
ECHO inriktar sig för närvarande på att tillhandahålla medicinsk utrustning och akut hälsovård , på stöd till inrättningar liksom vaccinering .
Insatserna inriktas dock alltmer på att upprätta ett självförsörjande hälsovårdssystem i provinsen .
UNMIK har redan tagit på sig en betydande roll på detta område .
Vidare har det i enlighet med återuppbyggnadsprogrammet inletts brådskande insatser på sjukhuset i Mitrovica i form av ett återuppbyggnadsprogram på 1 miljon euro .
Utvecklingen går långsamt på grund av de spända förbindelserna mellan de etniska grupperna i denna delade stad .
Kommissionen fortsätter dock sina insatser med stöd av UNMIK för detta projekt .
Vi hoppas att det en dag blir en symbol för att främja fördelarna med etnisk försoning .
Enligt europeiska gemenskapens uppskattning av skador uppgår de beräknade kostnaderna för återuppbyggnad av hälsovårdsinrättningar och anskaffning av utrustning till apotek och vårdcentraler till 4 miljoner euro .
Kommissionen skall nu inleda arbetet med biståndsprogrammen för år 2000 .
Vi tror att vi kan anslå en betydande summa till att förbättra hälsovårdssystemet .
Tonvikten kommer att ligga på långsiktiga reformer som täcker finansiering liksom utbildning och materialanskaffning inom hälsosektorn .
Arbete pågår redan tillsammans med UNMIK för att fastslå ett lämpligt bidrag från kommissionen för detta initiativ .
Herr kommissionär !
I morse framhöll ordförande Prodi bl.a. att vår förmåga till effektiva insatser sätts på prov på Balkan , att Europeiska unionens trovärdighet sätts på prov och att det är dags att låta ord och handling följas åt .
Vi har fått uppgifter om den höga spädbarnsdödligheten och barnadödligheten i Kosovo den högsta i Europa - men vi har också en allmän uppfattning om den humanitära katastrofsituationen i Kosovo .
Anser ni inte , herr kommissionär , att detta redan i sig allvarligt skadar vår trovärdighet och tilltron till vår förmåga att leva upp till våra löften ?
Och vidare , herr kommissionär , svarar den s.k. humanitära militära insatsstyrkan mot behoven i det katastrofdrabbade Kosovo ?
Anser ni att man kan rättfärdiga en så stor passivitet , när själva rätten till liv hotas på den europeiska kontinenten ?
Jag tror inte att vårt återuppbyggnadsorgan eller insatsstyrkan innan den , vilken har arbetat otroligt hårt i Kosovo , skulle anse det vara en riktig beskrivning av deras arbetsinsatser att antyda att de stått bredvid sysslolösa .
Jag är säker på att ärade ledamoten inte menade det .
Naturligtvis har hon helt rätt när hon säger att unionens trovärdighet står på spel med det som händer inte bara i Kosovo utan på hela Balkan .
Jag är mycket angelägen om att den hjälp vi tillhandahåller anländer snabbt och på ett sätt som ytterligare ökar våra hjälpinsatser .
Jag vill endast ta upp två punkter om situationen i Kosovo som vi håller på att försöka lösa så positivt som vi kan i överensstämmelse med WHO .
För det första är jag säker på att ärade ledamoten känner till att under 1990-talet underfinansierade regeringen i Belgrad hälsovårdssystemet i Kosovo och många albaner upptäckte att de inte fick någon hälsovård alls .
Till följd av detta inrättades ett parallellt hälsovårdssystem genom Moder Teresa organisationen .
Vad det således handlar om är inte bara följderna av konflikt utan resultaten av år av misskötsel och ständigt för litet investeringar .
Vidare , och jag är säker på att den ärade ledamoten känner till detta likaså , har några av de tragiska historier som man hört från Kosovo under de senaste veckorna inte handlat om barndödlighet under graviditet utan barndödlighet efter det att ett friskt barn fötts .
Detta gällde fall där kvinnor före eller under fientligheterna tragiskt dödade sina egna barn .
Vi har att göra med en fasansfull historia i Kosovo .
Vi måste arbeta så bra vi kan på hälsovårdsområdet och andra områden för att återställa något som liknar civila normer och civilt uppträdande , men det kommer inte att bli lätt .
Herr kommissionär !
Jag tackar er för ert svar på den första frågan från min kollega och även på den kompletterande frågan .
Jag har dock en del kontakter i Kosova och där säger man att de matpaket som delas ut bland annat av ECHO ofta är av undermålig kvalitet .
I vissa fall har man också hittat insekter och så i maten .
Känner ni till det ?
Är ni beredd att göra något åt det ?
Det är min första kompletterande fråga .
Min andra fråga gäller er hänvisning till återuppbyggnaden av sjukhuset i Mitrovica .
Ni känner kanske till att det sjukhuset ligger i den norra delen av staden och att , med tanke på det spända läget , Kosovoalbanerna inte alls får komma in där .
Vad gör kommissionen för att se till att även kosovoalbaner får tillgång till sjukhus ?
Som svar på den första frågan kommer jag själv att resa till Kosovo i början av nästa månad för ett andra besök och jag skall naturligtvis undersöka anklagelsen från ärade ledamoten om ECHO : s matpaket .
Jag har inte hört detta antydas förut , men det är en viktig punkt och jag skall naturligtvis undersöka den när jag är där .
Vidare förstår jag inte exakt vad ärade ledamoten menar om Mitrovica .
Jag var i Mitrovica för några månader sedan och såg själv situationen där .
Jag förde diskussioner med kommunala ledare från båda sidor , däribland ledaren för den albanska sidan som själv tidigare varit doktor och som var allmänt erkänd för det läkarjobb han hade utfört under fientligheterna och senare .
Så jag känner till de mycket allvarliga problem som finns på det sjukhuset och jag kan försäkra den ärade ledamoten att vi kommer att göra allt vi kan för att tillräckliga hälsovårdsinrättningar finns för alla i Kosovo , oavsett etnisk grupptillhörighet .
De speciella svårigheterna i Mitrovica , exempelvis albanska patienter som har problem att få komma till sjukhus , albansk personal har svårt att få arbeta där - är särskilt akuta problem .
Vi skall försöka lösa dem men det är inte lätt .
Fråga nr 37 från ( H-0029 / 00 ) : Angående : Turkiets blockad mot Armenien Genom avtalet om partnerskap och samarbete , som undertecknades den 12 oktober 1999 , främjar Europeiska unionen aktivt de sociala , ekonomiska och politiska förbindelserna med Armenien .
Vad gör kommissionen för att den turkiska regeringen skall häva den ekonomiska blockaden mot Armenien ?
Kommissionen stöder varje insats som syftar till att lösa konflikten mellan Turkiet och Armenien och beklagar att det fortfarande inte har skett någon normalisering av förbindelserna mellan dessa två länder .
Under rådande politiska förhållanden är det emellertid orealistiskt att tänka sig att gränsen mellan Armenien och Turkiet liksom den mellan Armenien och Azerbajdzjan kan öppnas utan en lösning på konflikten Nagorno-Karabach .
( PPE-DE ) .
( DE ) Herr talman !
Kommissionen skall ju också i framtiden föra förhandlingar på grund av anslutningen av Turkiet till Europeiska unionen .
Kommer den att sätta upp som villkor att diskussionen påbörjas först när blockaden här har avbrutits , ty när allt kommer omkring är vi alla grannar , och vi vill ju också vårda grannsämjan inom Europeiska unionen ?
Jag frågar alltså : Kommer kommissionen att göra detta till ett av villkoren för att förbättra de framtida samråden ?
Den viktigaste punkten är att stödja insatserna från OSSE : s grupp i Minsk för att hitta en lösning på Nagorno-Karabach konflikten och vi är beredda att hjälpa till på alla sätt vi kan .
Vi har även medverkat på ett omfattande sätt med utvecklingsstöd till Armenien inom ramen för Tacis-programmet .
Låt mitt svar speciellt sättas i samband med frågan om Turkiets anslutning till Europeiska unionen .
Situationen med Turkiets förbindelser med dess grannar kommer , såsom den ärade ledamoten begär , att noga granskas inom ramen för strategin för förberedelse för anslutning till unionen .
Såsom fastslås i Agenda 2000 - och jag citerar : " Utvidgning skall inte innebära att gränskonflikter förs in . "
Det uttalandet kan inte bli mer tydligt .
Men jag upprepar att det viktigaste bidraget vi kan göra är att försöka hjälpa till att lösa den konflikten som har orsakat sådana ekonomiska och humanitära skador .
Fråga nr 38 från ( H-0040 / 00 ) : Angående : Konsekvenserna av byggandet av Ilisudammen i Turkiet för de mänskliga rättigheterna Med tanke på att Turkiet nyligen gavs kandidatlandstatus , vad anser kommissionen om de konsekvenser som byggandet av Ilisudammen får för de mänskliga rättigheterna ?
Detta bygge kommer att medföra en stor omflyttning av den kurdiska befolkningen och av andra invånare i regionen .
Kommissionen har ingen information om effekten för befolkningen i regionen av att Ilisu- dammen byggs .
Vi skall dock överväga att ta upp frågan med de turkiska myndigheterna , tillsammans med andra frågor rörande regional utvecklingspolitik inom ramen för den nya strategin för Turkiets förberedelse för anslutning till unionen .
Jag har en närbesläktad punkt .
Den gäller dammens effekter för tillgång till färskvatten i regionen som helhet .
Som ni känner till kommer dammen att begränsa tillgången på vatten till Syrien och Irak i synnerhet .
Med hänsyn till hur ytterst instabil denna region är och många kommentatorers verkligt reella oro över att vi kommer att få se ett ökat antal konflikter , av så kallade " vattenkrig " , under de närmaste decennierna , vad anser kommissionen om den eventuella destabiliserande effekt både i Turkiet och i den bredare regionen som denna damm kommer att orsaka ?
Kan ni tala om ifall ni verkligen kommer att ta upp även denna fråga ?
Vi skall helt klart ta upp den punkt som den ärade ledamoten beskrivit .
Vi har fått höra oroliga frågor om detta och jag skall se till att den tas upp .
Det har också uttryckts betydande farhågor om den eventuella faran för de arkeologiska lämningarna i området .
Vi skall ta upp det också i de framställningar vi gör .
Ett antal andra vattenkraftsprojekt som planerats under de senaste 30 åren i Turkiet har framkallat oroliga frågor , som följderna för tvångsförflyttade bönder .
På det hela taget verkar dessa ha skötts relativt tillfredsställande och jag hoppas att samma sak kan gälla om detta projekt vilket - för att klargöra frågan - inte är ett projekt i vilket kommissionen deltar i någon form .
Vi tackar herr Patten för att han har företrätt kommissionen i besvarandet av dessa frågor .
Fråga nr 39 från ( H-0036 / 00 ) : Angående : Utkastet till en stadga om grundläggande rättigheter Det civila samhället ser med tillfredsställelse på utkastet till en stadga om grundläggande rättigheter och förhoppningen är att denna skall kunna anta de utmaningar som Europa kommer att ställas inför under det 2l : a århundradet .
Kan kommissionen mot denna bakgrund svara på följande frågor : Hur ser kommissionen på innehållet i stadgan ?
Vem skall stadgan gälla ?
Medborgare i Europeiska unionen eller i alla europeiska länder , med tanke på utvidgningen ?
Kommer den även att omfatta invandrare o.s.v. ?
Kommer stadgan att befästa Europeiska unionens sociala rättigheter eller kommer den att ha en bredare karaktär ?
Vilka mekanismer kommer att användas i stadgan för att tydligt säkerställa jämlikhet mellan de båda könen ?
Vad anser kommissionen om att införa stadgan i EU-fördraget ?
Liksom den ärade ledamoten , gläder sig kommissionen åt det beslut som fattats av stas- och regeringscheferna om att ta itu med utformningen av en EU-stadga om grundläggande fri- och rättigheter .
Stats- och regeringscheferna fastställde själva i Europeiska rådets slutsatser från Köln de stora linjerna för stadgans innehåll .
Enligt slutsatserna bör stadgan innehålla tre kategorier rättigheter : rätt till frihet , jämlikhet och rättslig prövning i enlighet med Europeiska konventionen om mänskliga rättigheter , rättigheter förbehållna unionens medborgare och ekonomiska och sociala rättigheter i enlighet med Europeiska socialstadgan och i Gemenskapens stadga om grundläggande sociala rättigheter för arbetstagare eftersom de inte endast omfattar mål för unionens verksamhet .
Kommissionen anser att den konvention som är ansvarig för utarbetandet av stadgan om grundläggande rättigheter bör respektera det mandat som lämnades av Europeiska rådet i Köln .
Det betyder dock inte att konventionen bör begränsas till en stadgande roll att bara räkna upp befintliga rättigheter från olika källor .
Såsom jag redan fått tillfälle att säga inför parlamentet är kommissionen övertygad om att konventionen i förekommande fall bör kunna anpassa och utveckla dessa rättigheter genom att ta hänsyn till aktuella omständigheter , i synnerhet tekniska och sociala förändringar .
Mot bakgrund av mandatet och det slutliga syftet med den text som skall läggas fram för stats- och regeringscheferna bör denna befogenhet utövas med försiktighet och från fall till fall .
De rättigheter som ges i stadgan kommer att tjäna åtminstone två kategorier .
Vissa rättigheter kommer att tillämpas för samtliga personer som befinner sig på unionens territorium , andra rättigheter kommer att kunna tillämpas endast för EU-medborgare .
Man skulle också kunna tänka sig att vissa ekonomiska och sociala rättigheter bara garanteras åt EU-medborgare och medborgare från tredje land som uppfyller vissa villkor .
Det är inte möjligt att på detta första stadium av utarbetandet av stadgan på förhand bedöma dess innehåll mer detaljerat .
Man kan dock påstå att bland annat principen om lika möjligheter och lika behandling av män och kvinnor säkert kommer att ingå i de rättigheter som skall garanteras av den framtida stadgan om grundläggande rättigheter i EU eftersom den redan finns bland de rättigheter , som garanteras i Fördraget om Europeiska gemenskapen och tillhörande rätt , och den utgör utan tvivel en gemensam konstitutionell tradition i medlemsstaterna .
Jag har redan sagt det också inför parlamentet att kommissionen är positiv till att stadgan skrivs in i fördraget .
Kommissionen är dock fullt medveten om att det slutliga beslutet i frågan åligger stats- och regeringscheferna .
Den svåra uppgift som konventionen har består således i att utarbeta en ambitiös och politiskt betydelsefull text , som direkt kan införlivas i fördragen .
I sitt yttrande om att samla en regeringskonferens i syfte att ändra fördragen påminner kommissionen om att Europeiska rådet skall uttala sig under år 2000 om införandet av vissa frågor i regeringskonferensens tidsplan , i synnerhet Europeiska unionens stadga om grundläggande rättigheter .
( Applåder ) Herr kommissionär !
Det är mycket betydelsefullt så här i början av det nya århundradet att Europas medborgare , män och kvinnor , uppmanas att ännu en gång definiera sina rättigheter och skyldigheter .
Jag hoppas verkligen att detta beslut från rådsmötet i Köln skall kunna genomföras .
Både globaliseringen och utvidgningen framtvingar en definition av dessa rättigheter .
Seattle innebär en verklig källa till problem i detta avseende , och jag hoppas att Europeiska rådets möte i Nice inte skall innebära ännu ett förlorat tillfälle .
För att medborgarna skall bli delaktiga i denna nya planering , skulle jag vilja veta vad de europeiska organen - närmare bestämt Europeiska kommissionen - har för förslag till social och ekonomisk modell för Europa under det 21 : a århundradet .
Jag har hört era allmänna riktlinjer , och jag skulle vilja fråga er vilken plats barnen , som självständiga individer , har i Europeiska kommissionens planering för den nya sociala modellen under det 21 : a århundradet .
Herr talman , fru ledamot !
Jag bör säga er mycket tydligt att , enligt min åsikt och såsom ordförande Prodi sade i morse , är utarbetandet av stadgan en politiskt mycket betydelsefull uppgift eftersom den visar att unionen placerar medborgarnas grundläggande rättigheter längst fram bland de politiska angelägenheterna för vårt gemensamma projekts framtid .
Inom den ramen måste man klart och tydligt säga på vilka kriterier man grundar sig för att välja rättigheter .
Jag tror att det väsentliga kriteriet är medborgarnas rättigheter gentemot de europeiska institutionerna .
Det är medborgarnas rättigheter såsom de anges i det europeiska projektet som fastställs i unionens fördrag .
Jag förstår er omsorg om barnens rättigheter .
Jag tror att flera delar av vårt arbete och framför allt av mitt arbete i egenskap av ansvarig för sektorn för rättsliga och inrikes frågor består i att se till barnens rättigheter .
Här kommer vi in på ett område där subsidiaritetsprincipen tillämpas fullt ut .
Varje medlemsstat har huvudansvaret för att fastställa sitt ansvar gentemot barnen .
När det gäller unionens ansvar som sådant tror jag att barnens rättigheter bör erkännas i stadgan genom att de områden beaktas där unionen kan tillföra ett mervärde till främjandet av den sociala , ekonomiska och till och med , i vidaste mening , medborgerliga situationen för barnen .
Jag hoppas att vi kommer att lyckas att anta den utmaning som ledamoten har ställt på kommissionen och på hela konventionen . Herr talman !
Jag har haft nöjet att höra kommissionären uttala sig ett antal gånger i denna fråga och jag håller mycket med honom och hans inställning .
Jag vill dock ställa en något annorlunda fråga .
Vi har just hört kommissionär Barnier säga att han är angelägen om att kommunicera bättre med människorna och att inrikta kommissionens informationspolitik mot de större frågor som gemenskapen arbetar med i år .
Skulle kommissionären anföra skäl för att någon del av kommissionens informationsbudget används för att informera och samråda med medborgarna i denna fråga om en medborgarstadga ?
Det är viktigt att människorna känner sig delaktiga i denna process .
Jag vet att själva konventet kommer att bidra mycket på detta område men den har inte de resurser som kommissionen har .
Kommer kommissionen att överväga att använda sin informationsbudget för att se till att människor blir intresserade av denna debatt ?
Det är kommissionens policy att främja en öppen och bred debatt om stadgan om grundläggande rättigheter , inte bara med icke-statliga organisationer utan också med medborgarna i ett projekt som är så omfattande som stadgan är .
Jag kan försäkra er att kommissionen kommer att göra sitt yttersta för att främja debatten om den framtida stadgan om grundläggande rättigheter .
Vi kan uppnå det bästa från båda världar genom att få en tydlig text och samtidigt en text som kan användas som ett rättsligt instrument .
Det finns ingen motsägelse mellan de två .
Vår utmaning är att sammanföra dem i den slutgiltiga versionen av stadgan .
Jag är mycket glad att veta att jag kan räkna med ert stöd i denna fråga .
Fråga nr 40 från ( H-0095 / 00 ) : Angående : Artiklarna 6.1 , 7.1 och 7.2 i Fördraget om Europeiska unionen I artikel 6.1 i fördraget står det att unionen bygger på principerna om frihet , demokrati och respekt för de mänskliga rättigheterna och de grundläggande friheterna .
Av de uttalanden som under de senaste åren gjorts av Jörg Haider och Frihetspartiet framgår det klart att dessa inte respekterar mänskliga rättigheter eller grundläggande friheter för tredjelandsmedborgare och minoritetsgrupper som är bosatta i Österrike .
Kan kommissionen därför ge besked om när kommissionen tänker åberopa artikel 7.1 om att " en medlemsstat allvarligt och ihållande åsidosätter principer som anges i artikel 6.1 " och yrka på att rådet med kvalificerad majoritet skall fatta beslut om att tillfälligt upphäva vissa av de rättigheter som Österrike har till följd av tillämpningen av detta fördrag , inbegripet rösträtten i rådet för företrädaren för Österrike ?
Herr talman , ärade kollegor !
Låt mig börja med att påminna er om kommissionens ståndpunkt när det gäller den nya österrikiska regeringen där ministrar från Jörg Haiders liberala parti ingår , något som upprepades i morse av ordförande Prodi .
Jag syftar givetvis på kommissionens uttalande från den 1 februari 2000 och vars huvudpunkter jag vill börja med att påminna om .
Kommissionen försäkrade på nytt och försäkrar i dag igen att man delar den underliggande oron i det portugisiska ordförandeskapets uttalande från den 31 januari .
Oron är berättigad och skälig .
Vi behöver inte påminnas om Jörg Haiders politiska bana och hans otaliga offentliga uttalanden , främlingsfientliga och rasistiska , med andra ord antieuropeiska .
Att ett klart extremistiskt , rasistiskt och främlingsfientligt parti kan komma till makten i en av Europeiska unionens medlemsstater är något som de övriga deltagarna i det europeiska projektet inte kan sluta att oroa sig över , på samma sätt som det inte är likgiltigt för Europeiska kommissionen .
För det andra så upprepade kommissionen , och upprepar igen , sitt åtagande att fortsätta fullgöra sina skyldigheter som fördragens väktare , särskilt det som åsyftas i artikel 6 och 7 i EU-fördraget .
En av de viktigare reformerna i Amsterdamfördraget var just de grundläggande principernas tydlighet , vilket är medlemsländernas gemensamma arv och institution för den kontrollapparat som krävs för att se till att de åtföljs och att en reaktion sker om någon av principerna kränks .
Kommissionen visade därmed i praktiken sin tillgivenhet för en av de grundläggande principerna : rättsstatens .
En sådan princip ålägger kommissionen att hålla sig inom de gränser som fastställts genom fördragen och det är i det här sambandet som uttalandet från den 1 februari skall ses .
Kommissionen är inte en stat , den varken kan eller bör agera som om den vore det .
Men för att besvara ledamotens fråga vill jag påminna om att den mekanism som instiftats i artikel 7.1 i EU-fördraget för att aktiveras kräver en bekräftelse på , jag citerar , " att en medlemsstat allvarligt och ihållande åsidosätter principer i artikel 6 " .
Jag upprepar , ett allvarligt och ihållande åsidosättande är ett oumbärligt villkor för att kommissionen skall kunna uppmana rådet att vidtaga åtgärder mot ett medlemsland .
För mig är det uppenbart att villkoren inte är uppfyllda för att tillämpa dem på situationen i Österrike .
Jag tror inte att jag misstar mig när jag säger att vi alla hoppas att ett sådant allvarligt och ihållande åsidosättande av de mänskliga rättigheterna och demokratin aldrig någonsin kommer att inträffa , varken i samband med Österrike eller något annat land inom unionen .
Jag vill dock försäkra er alla här i dag att min personliga ambition och kommissionens , som ordförande Prodi bekräftade i morse , är att göra allt som står i vår makt för att det inte skall bli nödvändigt att tillämpa artikel 7 .
Jag vill emellertid också säga att vi inte kommer att tveka att använda den om det behövs .
De värden som står på spel är alldeles för viktiga och grundläggande för att visa hänsyn eller kompromissa . § § Människor och regeringar bör värderas mera efter vad de gör än vad de säger .
I fallet med Österrike är uttalandena åtminstone motsägelsefulla .
Å ena sidan kan vem som helst av oss samla ihop ett antal upproriska meningar från det österrikiska liberala partiet .
Å andra sidan upprepar den nya österrikiska regeringen i sitt program sin ambition att försvara demokratin och de mänskliga rättigheterna .
Inom kort får vi ett ypperligt tillfälle att se vilken av de här två sidorna som är den rätta .
Jag tänker här på vilken ståndpunkt den österrikiska regeringen kommer att inta i rådet beträffande kommissionens förslag om ett åtgärdsprogram för kampen mot diskriminering samt två direktiv .
Ett som tillämpar principen om alla människors rätt till lika bemötande oavsett ras eller etniskt ursprung och ett annat som erbjuder ett skydd mot diskriminering vid anställning på grund av ras eller etniskt ursprung , religion och sexuell inriktning .
Det är relevanta dokument som godkänts i enlighet med artikel 13 i fördraget och där gemenskapen ges fullmakt att bekämpa diskriminering grundad på ras , etniskt ursprung , kön osv .
Låt mig avslutningsvis försäkra ledamoten om att kommissionen kommer att fortsätta att vara vaksam och vi kommer inte att sluta fullgöra våra skyldigheter , om detta skulle visa sig vara nödvändigt .
Jag tackar kommissionären för hans svar på min fråga .
Men är kommissionär Vitorino medveten om inte bara Haiders och Frihetspartiets uttalanden utan också deras gärningar ?
Haider har i själva verket varit verksam i ledningen i den södra provinsen Kärnten där han har lett en rasistisk och främlingsfientlig kampanj mot den slovensktalande minoriteten i den regionen som är österrikiska medborgare , där han har försökt att avskaffa tvåspråksutbildningen och där det har det skett en klar diskriminering mot romerbefolkningen och immigrantbefolkningen .
Kan kommissionären besvara två frågor .
För det första talade han om bekräftelse .
Kan han tala om hur den bekräftelsen skall ske och vem som skall göra den ?
För det andra , håller han inte med om att ifall den nuvarande regeringen på nationell nivå skulle bedriva den slags politik som Haider och Frihetspartiet bedrivit på regional nivå det klart skulle strida mot artikel 6.1 i fördraget i fråga om grundläggande fri- och rättigheter och det skulle falla på kommissionen att vidta nödvändiga åtgärder ?
Vi talar inte om uttalanden här .
Vi talar om gärningar av Frihetspartiet och Haider .
Jag anser det helt klart att det är kommissionens ansvar att noggrant följa utvecklingen av situationen i medlemsstaterna i enlighet med de förfaranden och normer som inryms i artikel 6 och som berättigar tillämpning av artikel 7 i fördraget .
Därför är jag helt förvissad om att kommissionen mycket noga kommer att kunna följa utvecklingen av situation i Österrike liksom i många andra medlemsstater .
Om något konkret fall av ständig kränkning av de mänskliga rättigheterna begåtts av regeringen i en medlemsstat kommer vi att var helt i stånd att reagera och agera därefter .
Jag förlitar mig inte bara på samarbetet från Europaparlamentets ledamöter utan även på samarbetet från icke-statliga organisationer som alltid har lämnat ett viktigt bidrag till kommissionens politik mot diskriminering .
Beträffande situationen i Kärnten , måste vi undersöka den närmare .
Ärade ledamoten tog upp frågan .
Skyddet för etniska minoriteter och för minoriteter som talar en särskilt språk är ett del av programmet och i de två direktiv som kommissionen har lagt fram för rådet .
Vi bör inte enbart inrikta denna debatt på den österrikiska frågan .
Den frågan kräver eftertanke , debatt och om så krävs , åtgärd .
Jag hoppas uppriktigt att alla medlemsstater skall ta möjligheten i fråga om denna handlingsplan och dessa två direktiv som kommissionen lagt fram för rådet att upprepa i klara och konkreta termer deras godkännande av handlingsplanen och direktiven och deras åtagande att bekämpa diskriminering , rasism och främlingsfientlighet varhelst det kan tänkas ske .
Tack så mycket , herr Vitorino , för ert värdefulla bidrag till frågestunden .
Andra delen Frågor till Wallström Fråga nr 41 från ( H-0021 / 00 ) : Angående : Elektriskt och elektroniskt avfall För varje år som går står EU inför en allt större mängd elektriskt och elektroniskt avfall ( 6 miljoner ton 1998 ) som framför allt beror på apparaterna blivit föråldrade i allt snabbare takt .
Miljöproblemen till följd av att dessa apparater förbränns eller slängs på soptippen beror i främsta rummet på att de innehåller farliga ämnen ( bly , kadmium , kvicksilver , hexavalent krom , PVC och halogenerade flamskyddsmedel ) .
Ett utkast till förslag till direktiv i syfte att reglera administrationen av dessa avfall gav upphov till tre på varandra följande versioner , den senaste från juli 1999 .
Kan kommissionen förklara varför administrationen av det här projektet tagit så tid , trots att det i princip borde ha varit klart 1998 ?
Stämmer det att den amerikanska regeringen motsätter sig de flesta bestämmelser i det nuvarande förslaget och att den till och med hotar att dra EU inför WTO ( för brott mot artikel XI i GATT-avtalet och artikel 2.2 i avtalet om tekniska handelshinder ) ifall förslaget antas ?
Kommissionen håller med parlamentsledamoten om att den nuvarande hanteringen av elektriskt och elektroniskt avfall inom Europeiska unionen orsakar betydande miljöproblem .
Kommissionen har därför beslutat att utarbeta ett förslag i ämnet och har sedan 1997 tagit upp frågan med alla berörda parter .
Resultaten från denna debatt och de grundliga efterforskningar som görs på området granskas nu av kommissionen .
Vissa delar av förslaget har utsatts för kritik , bland annat utfasningen av vissa tungmetaller och bromerade flamskyddsmedel samt tillämpningen av principen om tillverkarens ansvar för hanteringen av elektriskt och elektroniskt avfall .
Förenta staternas delegation vid Europeiska unionen har ställt sig tveksam till några punkter i det senaste samrådsdokumentet , bland annat just utfasningen av ovannämnda ämnen och vissa frågor som gäller principen om tillverkarens ansvar .
Förenta staternas huvudargument i detta sammanhang är att de ifrågavarande bestämmelserna påstås vara oförenliga med internationell handelsrätt .
Kommissionen har för närvarande delegationens argument under övervägande .
Låt mig tillägga att mina planer är att före påsk för kommissionen kunna presentera ett förslag om hantering av elektriskt och elektroniskt avfall .
Min fråga gällde just den amerikanska regeringens reaktion på texten i det förberedande projektet .
Det finns nämligen tre förberedande texter och den sista enligt min vetskap från juli 1999 .
Är det således denna text som ni skall lägga fram eller en ändring i förhållande till den ursprungliga versionen ? .
Den tredje versionen var nämligen redan svagare än den andra versionen till följd av den amerikanska industrins anmärkningar , som följdes upp av den amerikanska regeringen .
Jag vill i synnerhet påpeka att , när ni talar om den internationella rätt med vilken det sägs att texten inte överensstämmer , syftar ni nämligen på Världshandelsorganisationens regler .
Den amerikanska regeringens påståenden gäller det faktum att det skulle vara att gå emot WTO : s regler att på sikt förbjuda förekomsten av farliga ämnen i elektriskt och elektroniskt avfall .
Det bekymrar mig personligen eftersom det skulle betyda att om man antar en text står man ständigt under hot om en attack inför Världshandelsorganisationen , och det försvagar således fullständigt den europeiska miljölagstiftningen , i synnerhet detta förslag .
Tack för följdfrågan .
Det är viktigt att jag får tillfälle att svara på den .
Det är klart att i en process som denna , där vi diskuterar en mycket stor avfallsström i Europa av både elektriskt och elektroniskt avfall , pågår en ständig dialog mellan olika inblandade parter .
Vi har haft en bra dialog och har utvecklat ett förslag under processens gång .
Vissa avsnitt har stärkts , andra har vi kanske fått kompromissa litet för mycket med .
Vi håller fortfarande på att skriva på texterna , och dialogen med de olika inblandade parterna pågår ända in i sista minuten .
Jag vill säga att jag inte anser att Förenta staternas inblandning i denna fråga skall låta oss styras på ett sådant sätt att vi inte tar tillräcklig miljöhänsyn .
Jag värjer mig verkligen mot att man ständigt skall kunna hänvisa till WTO och handelsregler för att förhindra att vi i EU skaffar oss radikala miljöbestämmelser .
Min utgångspunkt är att vi skall göra det .
Jag är emellertid beredd att lyssna på alla argument .
Jag har exempelvis nyligen träffat företrädare för elektronikbranschen .
De lämnade förslag - också praktiska - till hur man skulle kunna förbättra vårt förslag .
Jag vill dock bestämt tillbakavisa påståendet att jag skulle låta Förenta staterna styra utformningen av vårt direktiv .
Det är faktiskt så att jag menar att vi måste visa vägen , vilket också kommer att prägla det slutgiltiga förslaget .
Fråga nr 42 från ( H-0026 / 00 ) : Angående : Gender och miljö Så gott som samtliga aktörer i Rio- och Kyotoprocesserna - enskilda organisationer , medborgarrörelser , regeringar Världsbanken , FN och hjälporganisationer - ansåg att kvinnor i högre grad skall delta i beslutsfattande inom miljöområdet.Fler kvinnor i beslutsfattande positioner inom olika miljöorgan gör att de förhärskande manliga referensramarna utvidgas till att omfatta inte bara frågor som berör företagande utan även sociala rättvisefrågor .
Är kommissionen beredd att anta en handlingsplan för att öka kvinnors aktiva deltagande i beslutsfattande även inom miljöområdet .
Kommissionen har sedan 1988 ett handlingsprogram för lika möjligheter för kvinnor och män .
Med hjälp av det nuvarande programmet , som omfattar åren 1997 till 2000 , försöker man utveckla en arbetskultur , som innebär att både manliga och kvinnliga värden integreras , och att hänsyn tas till könsspecifika behov .
Ett av programmets syften är att utarbeta och övervaka metoder , strategier och åtgärder , som främjar en jämn könsfördelning i beslutsprocessen , däribland på högre befattningar .
Inom ramen för detta handlingsprogram utarbetar varje enskilt generaldirektorat en särskild åtgärdsplan .
Ett av målen i åtgärdsplanen är att öka antalet kvinnor i ledande ställning .
Den nya kommissionen har som mål att fördubbla antalet kvinnliga chefer under sin mandatperiod .
Denna linje drivs särskilt aktivt på generaldirektoratet för miljö , där för närvarande 60 procent av direktörerna och 20 procent av enhetscheferna är kvinnor .
Vår politik är att gynna rekryteringen av kvinnor till administrativa tjänster för att skapa en reserv av lämpliga kandidater för framtida chefstjänster .
För närvarande är 24,5 procent av våra A-tjänstemän kvinnor .
Vi hoppas att antalet kommer att öka stadigt .
Vi anstränger oss dessutom för att locka kvalificerade kvinnor att delta i de samrådsforum som vi organiserar .
När det gäller våra externa partners kan vi bara föregå med gott exempel och uppmuntra deras ansträngningar att demokratisera sina beslutsprocesser .
När det gäller mer allmänna frågor om integrering av jämställdhetsperspektivet , känner ni säkert till att denna princip ingår i Amsterdamfördraget .
I artikel 3 i fördraget anges att gemenskapen i all verksamhet som avses i denna artikel skall syfta till att undanröja bristande jämställdhet mellan kvinnor och män och att främja jämställdhet mellan dem .
Kommissionen ger sitt fulla stöd till ansträngningarna på detta område och håller på att undersöka om specifika åtgärder kan vidtas på miljöområdet .
Naturligtvis vill jag passa på att säga att jag uppskattar den roll som Europaparlamentets kvinnoutskott , och inte minst dess ordförande , spelar .
Låt mig bara påminna om att när den nuvarande kommissionen så småningom godkändes fick varje kommissionär en fråga från kvinnoutskottet om hur de inom just sitt verksamhetsområde skulle sköta jämställdheten .
Vi kommer noggrant att granska varje kommissionär , så jag vill härmed förvarna även de andra kommissionärerna .
Tack så mycket för svaret !
Jag tolkar det faktiskt som ett ja till att det är en handlingsplan som behövs - en handlingsplan för att få fler kvinnor att delta inom specifika miljöområden .
Låt mig också säga att Pekingdeklarationen understryker vikten av att ha institutionell kapacitet för att ta med ett jämställdhetsperspektiv i all miljöprogrammering .
Miljöinstitutioner saknar ofta kunskaper och procedurer för att inkorporera ett sådant perspektiv i sitt dagliga arbete .
Jag vill naturligtvis veta om kommissionären är villig att integrera jämställdhetstänkandet i miljöpolitiken och i miljöprogrammen .
Detta är viktigt .
Om hela politiken skall genomsyras , tror jag att det är särskilt viktigt att cheferna på hög nivå har denna grundläggande kunskap . .
Naturligtvis är min bild av mainstreaming att detta måste prägla allt vi gör .
I den plan som utarbetas på mitt generaldirektorat spelar jämställdhetsfrågorna en mycket viktig roll .
Jag är också beredd att själv gå in och exempelvis leda seminarier i ledarskap eller andra ämnen för att uppmuntra kvinnor att ta på sig vidare uppgifter inom kommissionen .
Om vi skall kunna motivera alla , tror jag att det är väldigt viktigt att detta budskap sänds hela vägen uppifrån och ned - eller nedifrån och upp om du så vill .
Min bild av miljöarbete i stort är att det många gånger domineras av kvinnor .
Det handlar om att detta måste fortplantas , så att kvinnor har en chans att också få chefsjobb eller komma till högre positioner inom miljöarbetet .
Jag vill påstå att vår åtgärdsplan avspeglar detta , men den kan säkert göras bättre .
Jag har en viss erfarenhet av att upprätta planer och följa upp dem .
Jag hoppas att detta skall komma till nytta .
Fråga nr 43 från ( H-0045 / 00 ) : Angående : Området vid mynningen av floden Boyne och företaget Drogheda Området vid mynningen av floden Boyne är klassificerat som ett särskilt skyddsområde enligt direktivet om vilda fåglar och man överväger för närvarande att klassificera det som ett särskilt bevarandeområde enligt habitatdirektivet på grund av dess internationella betydelse .
Marindepartementet , grevskapsrådet i Louth och företaget Drogheda har godkänt uppförandet av en ny hamn i det särskilda skyddsområdet och till och med avskaffandet av en strandremsa i Stegrennan , som nyligen införlivades i det särskilda skyddsområdet på kommissionens uttryckliga uppmaning .
Dessutom har man uppfört ett mycket stort lagerhus .
Det har visat sig vara svårt att få tag på byggnadstillståndet för detta lager , och Drogheda planerar samtidigt annan infrastruktur .
Hur kan kommissionen säkerställa att sådana projekt som finansieras via strukturfonderna inte går stick i stäv mot miljöskyddsbehoven i området ?
Är kommissionen beredd att inställa finansieringen helt och hållet i väntan på att utvecklingsplanerna för detta område skall ses över ?
Kommissionen känner till uppförandet av hamnen , men vet inget om det lagerhus , eller den övriga infrastruktur som parlamentsledamoten nämner .
Hamnens uppförande får stöd från strukturfonderna och medför i huvudsak att utloppet i floden Boynes mynning muddras och att muddermassorna mellanlagras på Stegrennans strandremsa .
Floden Boynes mynningsområde är klassificerat som särskilt skyddsområde enligt direktivet om vilda fåglar .
Detta innebär att man vid all exploatering i eller vid Boynesmynningen , som kan komma att påverka det särskilda skyddsområdet , måste beakta de skyddsbestämmelser för området som fastställts i gemenskapens habitatdirektiv .
Sedan 1998 har det till kommissionen kommit in ett antal klagomål , där man hävdar att hamnanläggningen kommer att skada Stegrennans strandremsa , som numera ingår i det särskilda skyddsområdet , och att man inte har beaktat de relevanta skyddsbestämmelserna .
Efter att ha granskat dessa klagomål under 1998 och i början av förra året - projektet erhöll under denna tiden inga medel från strukturfonderna- blev kommissionen på sommaren 1999 övertygad om att man vid uppförandet av hamnen hade beaktat de relevanta skyddsbestämmelserna .
En detaljerad miljökonsekvensbedömning hade gjorts .
Den mest negativa följden av projektet , förlusten av Stegrennans strandremsa , skall endast vara tillfällig , och entreprenören är skyldig att helt återställa strandremsan .
På kommissionens uppmaning införlivades Stegrennansstrandremsa formellt i Boynesmynningens särskilda skyddsområde , från vilken den tidigare hade varit utesluten .
För att uppväga de negativa effekterna av strandremsans tillfälliga försvinnande på berörda fågelpopulationer var det dessutom meningen att andra livsmiljöer i mynningsområdet skulle förbättras .
Sedan sommaren förra året har emellertid den sistnämnda åtgärden varit omtvistad .
Först drog de irländska myndigheterna tillbaka sitt tidigare förbättringsåtagande .
De förnyade sedan sitt åtagande efter det att en icke-statligt irländsk miljöorganisation hade anfört klagomål inför irländsk domstol .
Det nya åtagandet innehöll dock smärre ändringar , som i sin tur ledde till ytterligare ett klagomål .
Mot bakgrund av att Irland har åtagit sig att vidta kompensationsåtgärder , och med tanke på att andra frågor redan har lösts , vill kommissionen för närvarande inte föreslå att man ställer in finansieringen från strukturfonderna .
Kommissionen vill dock reda ut spörsmålet om kompensationsåtgärden avseende förbättrade livsmiljöer med de irländska myndigheterna , särskilt i ljuset av den ännu oavslutade processen inför irländsk domstol .
Jag förstår inte riktigt det som kommissionären sade .
Den gyttjiga strandremsan vid Stregrennan , som gjordes till ett särskilt skyddsområde på kommissionens begäran har förstörts helt i detta skede .
Det är uppenbart att de aktiviteter som har skett där klart bryter mot EG-direktiven .
Ni säger att det inte kommer att anslås mer medel .
Jag skulle vilja veta om ni tänker stoppa finansieringen helt i detta skede tills det blir en ordentlig utredning .
Om inte , varför inte ?
Om ni tänker göra det , när exakt kommer ni att göra det ?
Är det rätt och lämpligt att det departement som äger företaget också är den myndighet som utfärdar tillståndet och även den myndighet som praktiskt taget tar emot pengarna från EU och ger det till ett företag som det äger till 100 procent ?
Är detta rätt och lämpligt ?
Vad anser ni om det ?
Varje bidrag från EU till projektet måste stoppas eftersom det klart bryter mot EG-direktiven .
Även det område som utsetts som särskilt skyddsområde av kommissionärerna har förstörts .
Skadestånd efteråt kan inte gottgöra den skada som uppstått .
Den första rättsliga utmaningen kom efter det att arbetet med att uppföra hamnen inletts tidigt på hösten 1999 utan att förbättringar i form av kompenserande livsmiljöer inrättats .
Till följd av det gick de irländska myndigheterna med på att på nytt börja avlägsna marskgräset men denna gång på mekanisk väg .
Användningen av mekaniska hjälpmedel ledde till ytterligare ett klagomål - det är vad jag tog upp även i mitt första svar - grundat på argumentet att man genom mekaniskt avlägsnande skulle skada underliggande gyttjemark och orsaka ekologiskt skadlig spridning av marskgräset i flodmynningen .
Det finns hittills inget slutgiltigt resultat på detta klagomål .
Beslut om nödvändiga kompensationsåtgärderna är en fråga för de nationella myndigheterna och kräver inget föregående godkännande av kommissionen .
Kommissionens roll är att se till att de normer som gäller enligt fågeldirektivet beaktas fullt ut och uppenbarligen skulle det bli problem med kompensationsåtgärder som i sig själva orsakar skada .
I detta fall föreslår kommissionen att få ytterligare klargöranden från de irländska myndigheterna om det aktuella läget med kompensationsåtgärderna och eventuella problem med det mekaniska avlägsnandet av marskgräs .
Vi är för närvarande inte beredda att föreslå att man ställer in finansieringen från strukturfonderna .
Herr talman !
Tyvärr är det speciella fall som McKenna tog upp inte ett isolerat sådant .
Det finns andra exempel på naturskydd på särskilda vetenskapliga områden där skador uppstått till följd av finansiering från EU .
Kommer kommissionen att överväga att utfärda föreskrifter till alla medlemsstater om att om den i framtiden upptäcker att man bryter mot de europeiska miljödirektiven eller tillämplig miljökonsekvensbedömning inte skett kommer den inte bara att inställa vidare finansiering utan även att upphäva beslut om redan beviljade medel , med andra ord , återkräva pengar från medlemsstaterna ?
Det är endast en sådan åtgärd som kommer att avskräcka denna praxis i framtiden . .
Detta är en mycket viktig fråga .
Som Europaparlamentarikerna säkert känner till , gick det under förra året ut ett gemensamt brev från våra föregångare i kommissionen , Ritt Bjerregaard och Monika Wulf-Mathies angående förhållandet mellan strukturfonderna , pengar från strukturfonderna och skyddet i habitat- och fågeldirektiven .
Det budskap som sändes ut i detta gemensamma brev gäller fortfarande .
Vi kan inte med ena handen dela ut pengar och med den andra dra länderna inför domstol och kanske så småningom få böter utdömda .
Det är därför viktigt att detta står i samklang .
Naturligtvis kan svåra avvägningsfall bli följden .
Som jag ser det , är dock den främsta effekten att länderna tänker sig noga för och framför allt ser till att skicka in sina listor över Natura 2000-platser , så att vi har möjlighet att övervaka och följa upp på ett ordentligt sätt .
Där brister Irland i likhet med andra medlemsländer , men vi hoppas att vi skall kunna se resultat av denna påtryckning .
Jag vill ännu en gång påpeka att det som stod i detta brev fortfarande är giltigt .
Det tillåter inte arbetsordningen .
Ni får lov att diskutera det utanför plenisalen , fru ledamot .
Frågor till Barnier Fråga nr 44 från ( H-0020 / 00 ) : Angående : Partnerskap och den tredje gemenskapsstödramen i Grekland Den nya förordningen ( EG ) 1260 / 1999om allmänna bestämmelser för strukturfonderna betonas , i motsats till i föregående förordning , att partnerskap skall förstärkas och att regionala , lokala och övriga behöriga offentliga myndigheter , arbetsmarknadens parter , näringslivets organisationer och alla andra relevanta organ skall delta i att förbereda och finansiera , övervaka och utvärdera stödåtgärder .
Enligt upprepade klagomål från lokala myndigheter är förfarandena vad gäller den nya grekiska gemenskapsstödramen dock oförändrade och " parternas " roll framhävs inte alls .
Kan kommissionen , mot denna bakgrund , svara på följande frågor : Har den grekiska regeringen tillfogat några ändringar till förfarandena för att bredda partnerskapens sammansättning så att dessa i synnerhet även omfattar lokala myndigheter och andra representativa organ ?
Vad innebär vidare de lokala myndigheternas ökade roll i förberedelsen och finansieringen av den tredje gemenskapsstödramen ?
Vilka åtgärder kommer slutligen kommissionen att vidta för att säkerställa ökat deltagande från " parternas " sida inom alla förfaranden som den nya gemenskapsstödramen omfattar ?
Tillåter ni mig att förlänga Margot Wallströms svar till ordförande David Martin med en mening för att säga att eftersom det handlade om en gemensam skrivelse mellan våra båda föregångare anser jag i egenskap av efterträdare till Wulf-Mathies att skrivelsen förvisso fortfarande är giltig och att jag i gott samförstånd skall ta itu med att tillsammans med Margot Wallström kontrollera om de projekt som finansieras genom strukturfonderna är förenliga med EU : s miljödirektiv och -politik .
Det är också en före detta miljöminister som svarar er , ordförande Martin .
Jag skulle nu bara vilja säga några ord till Alavanos som förlåter mig denna inträngning i ett annat ämne för att säga till svar på hans fråga att kommissionen inom ramen för förberedelsen av den nya programplaneringsperioden förvisso har sett till och kommer att se till att partnerskapsprincipen tillämpas .
Jag tillåter mig att här påminna om , men ni vet det , att anslutningen av de regionala och lokala myndigheterna till gemenskapens verksamhet utgör en av de främsta beståndsdelarna i den nya förordningen för strukturfonderna från Berlin .
När det mer speciellt rör tillämpningen av partnerskapsprincipen vad gäller den kommande gemenskapsstödramen i Grekland har kommissionen kunnat notera att de offentliga myndigheterna i stor utsträckning har fått bidra till utarbetandet av den grekiska planen för regional utveckling för perioden 2000-2006 .
Alavanos vet att jag för övrigt har varit där två gånger under ganska tragiska omständigheter till följd av jordbävningsdramat och under dessa besök har jag kunnat diskutera med den grekiska regeringen och påminna om angelägenheten att beakta partnerskapsmålet och -kravet .
När det gäller följande faser , herr ledamot , det vill säga utarbetandet av de nationella och regionala programmen räcker det inte att detta mål beaktas på nationell och teoretisk nivå , det måste göras konkret i de program som utgår från gemenskapsstödramen på de nationella , regionala och lokala planen .
När det gäller uppföljning och förvaltning av programmen har jag ännu inte i detta ögonblick mottagit de nationella bestämmelser som föreslagits av den grekiska regeringen för tillämpning av artikel 8 i den nya förordningen .
Jag kan meddela er att jag , inom ramen för förhandlingarna om den tredje gemenskapsstödramen som för närvarande pågår , har bett att bestämmelserna i samband med partnerskapsprincipen skall respekteras fullt ut , inbegripet för de regionala och lokala myndigheterna och inbegripet för allt som rör icke-statliga organisationer och sammanslutningar .
Denna princip bör sålunda överföras inom ramen för den tredje gemenskapsstödramen , i synnerhet genom deltagande av samtliga partner till uppföljningskommittén .
Herr ledamot , det är det svar jag kan ge er .
Jag tackar kommissionären .
Jag ifrågasätter inte alls hans avsikter och insatser som rört sig i en positiv riktning .
Men situationen är helt annorlunda .
Just nu får vi uppleva en stark maktkoncentration och både statlig och partipolitisk maktberusning när det gäller bidragen från Europeiska unionen .
Jag kan inte förmedla TV-programmen här , men jag har tagit med mig några grekiska tidningar till er från veckorna före valet .
I alla Greklands söndagstidningar kan man läsa : Ministeriet för offentliga anläggningsarbeten om strukturfonden : tack vare ministern ; Jordbruksministeriet : tack vare jordbruksministern - några veckor före valet - Telekommunikationsministeriet : tack vare telekommunikationsministern ; Utbildningsministeriet : tack vare utbildningsministern och så ett fotografi på ministern ; Arbetsmarknadsministeriet : tack vare arbetsmarknadsministern , ett fotografi på ministern och ett på biträdande ministern och bakom allt detta emblemet för gemenskapens strukturfonder .
Vi har bara några veckor kvar till valet .
Propaganda för parti och kandidater , som finansieras med hjälp av gemenskapens strukturfonder .
Jag ställer en fråga till kommissionären : Kommer kommissionen att tiga ?
Kommer kommissionen att ta upp det här med den grekiska regeringen , eller kommer denna kommission att utvecklas i samma patologiska riktning som den föregående ?
Herr Alavanos , jag har förstått att ni kastar de dokument åt vänster som ni har nämnt .
Det skulle vara mig ett nöje om vi ville ge mig dem så att jag kan läsa dem - ja , jag kommer att låta översätta dem - och att jag tittar på vad som liknar information , kommunikation , som jag bara kan glädja mig åt i egenskap av kommissionär med ansvar för regionalpolitik , och propaganda .
Och därefter om det är absolut nödvändigt att jag gör det kommer jag att lämna synpunkter eller rekommendationer till den grekiska regeringen .
Jag skulle således bli mycket lycklig , herr ledamot om ni kunde ge mig dokumenten eller också går jag och hämtar dem om en stund på golvet i er grupps rad .
Därmed sagt att jag trodde att er fråga mer avsåg partnerskapet .
Bortom dessa frågor förbundna med den förberedande valperioden som ni anger , säger jag än en gång att jag är bekymrad över att de regionala och lokala myndigheterna är anslutna på samma gång som icke-statliga organisationer .
Men jag kan inte heller skriva något annat än det som står i den allmänna förordningen om strukturfonderna och anger att kommissionen skall arbeta med medlemsstaternas regeringar och att det är den grekiska regeringen som jag har till partner , såsom första partner .
Sedan måste jag försäkra mig om att partnerskapet sprids , eftersom jag är decentraliserad skall jag försäkra mig om det .
Jag kan inte göra annat än att arbeta med den grekiska regeringen .
Jag tror att vår kollega Alavanos kommer att ge kommissionsledamoten alla dessa uppgifter , så att han kan ta ställning till dem , för det är faktiskt fråga om propaganda och inte något slags reklam för gemenskapens program .
Men i själva sakfrågan vill jag be kommissionären att ta hänsyn till följande : att Grekland i fråga om samtliga både nationella och regionala program betraktas som en enda region som - i partnerrelationen till Europeiska unionen ­ företräds av centralförvaltningen , av centralregeringen .
Detta innebär att varken de lokala självstyrelseorganen eller - än mindre - icke-statliga organisationer , som t.ex. de jordbrukskooperativa företag som skulle kunna vara intresserade av en utveckling av jordbrukssektorn , deltar i utarbetandet av förslag i fråga om gemenskapens tredje stödprogram och inte heller har medverkat i fråga om gemenskapens tidigare stödprogram .
Hur kan kommissionen hantera denna fråga ?
Än en gång Theonas , säger jag om vad jag sade till Alavanos , jag kommer att nära titta på och , om det behövs , kommer jag att inom ramen för och med iakttagande av strukturfondernas förordning lämna synpunkter på den användning man gör , inte av strukturfonderna som ännu inte har använts utan om förhandlingen före tilldelningen av dessa strukturfonder .
Men än en gång , jag måste respektera den nationella myndighet med vilken jag skall genomföra förhandlingen .
Jag kommer ändå att se det hela på ett objektivt sätt .
Herr Theonas , om ni har rekommendationer eller förslag om anslutning av den ena eller andra strukturen - ni talade om kooperativ om jag förstod rätt - är jag öppen och jag är beredd , på grundval av förslag från Europaparlamentets ledamöter , ni har er roll och jag har min , att ta över förslag så länge de respekterar tanke och innehåll i förordningen om strukturfonderna .
Varför skulle jag inte säga att vi från den grekiska regeringens sida tidigare år har noterat vissa brister när det gäller tillämpningen av den nya förordningen och den föregående förordningen om anslutning av företrädare för det civila samhället .
Jag säger det objektivt och när man upptäcker ett problem eller brister måste man avlägsna problemet eller bristerna .
Jag skall således se till att det blir gjort inom ramen för genomförandet av den nya gemenskapsstödramen .
Fråga nr 45 från ( H-0041 / 00 ) : Angående : Finansiering från strukturfonderna av forskning på kärnkraftsområdet Kan kommissionen bekräfta att det i den senaste programperioden för strukturfonderna , 1994-1999 , inte utgick något stöd till forskning inom kärnfusion och kärnfission ?
Kan den också vid de pågående förhandlingarna med medlemsstaterna om planer och program för den nya perioden , 2000-2006 , arbeta för att inte bevilja några finansieringsåtgärder för den här typen av forskning ?
Vilken roll kommer å andra sidan strukturfondsstödet att spela för att främja förnybara energikällor ?
Kan man förvänta sig att finansieringen från strukturfonderna inom energipolitiken inriktas på att främja regionala och förnybara energikällor ?
Kommer stöd från strukturfonderna även att utgå till de stora näten för energiöverföring ? ¿ Jag skulle vilja svara Isler Béguin på den första punkten och påminna henne om att förbättringen av den vetenskapliga grunden och regionernas tekniska kapacitet i syfte att öka konkurrensförmågan utgjorde en av gemenskapens prioriteringar under den föregående programplaneringsperioden .
Det stöd som tilldelas genom strukturfonderna till förmån för teknisk sammanhållning , det vill säga forskning och teknisk utveckling vad gäller gemenskapsstödramarna under denna period uppskattas till omkring 7,5 miljarder euro .
Det är ungefär 6 procent av det sammanlagda gemenskapsbidraget , fru ledamot .
Vad beträffar just ert bekymmer vill jag säga er att liksom under den föregående perioden har kommissionen inte för avsikt att direktfinansiera forskning och teknisk utveckling på området för fusion eller fission i samband med kärnkraft genom strukturfonderna .
Det fortsätter att vara på medlemsstaternas förvaltningsmyndigheters ansvar att välja de projekt som genomförs inom ramen för dessa gemenskapsstödramar .
Fru ledamot , även om det inte utgör en prioritering för gemenskapen kan en medlemsstat besluta att finansiera projekt för forskning och utveckling på den civila kärnkraftens område så länge som dessa projekt bidrar till den regionala utvecklingen och utan att för den skull systematiskt informera kommissionen om det .
När det gäller er andra punkt , som ni vet intresserar mig och fortsätter att intressera mig i hög grad , de förnybara energierna , läggs kommissionens tillnärmning fram i dokumentet om strukturfonderna och deras samordning med Sammanhållningsfonden .
De avser att investeringar inom sektorn för förnybara energier bör uppmuntras eftersom de främjar utveckling av lokala resurser där de bidrar till beroendeminskning i förhållande till energiimport och är också sysselsättningsskapande på lokal nivå .
Jag har kunnat kontrollera det , till exempel vid ett besök i Portugal för några dagar sedan på Azorerna , där det handlar om en naturlig källa till förnybar energi .
Strukturfondernas bidrag till förmån för en större genomträngning på marknaderna av förnybara energier , underströks också i kampanjen för säljstart för förnybara energikällor som inletts av generaldirektoratet för transport och energi .
När det slutligen gäller de stora energinäten , avses också i riktlinjerna ett finansiellt deltagande genom fonden för utveckling av transportnät för energi , när denna bidrar till att minska beroendet gentemot en extern leverantör eller för att bekämpa isoleringseffekter .
Det gäller i synnerhet för den region som jag nämnde , Azorerna , men också för samtliga områden i de yttersta randområdena och , jag vill tillägga , också för vissa regioner som är handikappade genom isolering på grund av berg , till exempel .
Herr kommissionär !
Jag har hört ert svar men , å andra sidan , om jag ställde frågan är det just för att vi är oroliga , eftersom ett projekt kallat " International Thermonuclear Experimental Reactor " förekommer inom ramen för betänkandet om den tredje gemenskapsstödramen för forskning .
Det uppgår till flera miljarder euro och områden som kan få strukturfonder , såsom mål 1-områdena , skulle kunna få ta emot denna typ av anläggning .
Det som vi skulle vilja veta , det är nämligen om kommissionen skulle vara beredd att finansiera denna typ av projekt inom ramen för anläggningen av denna forskningsplats och kanske inte direkt inom den specifika ramen för " kärnforskning " .
Herr Barnier , förlåt mig men ni svarade inte helt och hållet på den andra delen av min fråga om de stora transportnäten för energi .
Skulle ni kunna ge ett svar på detta ?
Ni oroar er över att få veta om vi skall finansiera en anläggning av kärnkraftverk någonstans med strukturfonder ?
Jag förenklar .
Man kan säga att det inte är fråga om det .
Jag har sagt er att projektvalet är medlemsstaternas sak utifrån förordningen om strukturfonderna .
Kommissionens enheter är följaktligen inte systematiskt informerade om samtliga valda projekt .
Ni gör dock rätt i att fråga mig , det är ert arbete och mitt är att svara .
Liksom det har skett i det förflutna , måste medlemsstaterna svara då kommissionen frågar dem eller begär klargöranden .
Jag skall således gå litet längre än det förtroende som vanligen delas mellan medlemsstaterna och kommissionen , och om den speciella punkt som ni nämner skall jag se efter exakt vad det handlar om .
Den medlemsstat eller de berörda medlemsstaterna måste då svara mig och jag kommer genast att hänvisa svaret till er .
Jag trodde mig ha svarat på frågan om de stora näten .
Energisituationen varierar kraftigt beroende på område i Europeiska unionen och stödet från fonderna skulle i vissa fall och för vissa områden kunna berättigas i synnerhet i de fall där anslutningen till de grundläggande energinäten ännu är underutvecklad .
Det är det svar jag kan ge om bandet mellan de stora näten och strukturfonderna .
Fråga nr 46 från ( H-0052 / 00 ) : Angående : Strukturfonderna och additionalitetsprincipen Mot bakgrund av kommissionens svar nyligen på min skriftliga fråga om strukturfonderna och additionalitetsprincipen undrar jag om kommissionen planerar att försöka ändra på reglerna om additionalitet .
Skulle kommissionen ställa sig positiv till ändringar i bestämmelserna för att se till att additionalitetsprincipen gäller inte bara på medlemsstatsnivå utan även inom medlemsstater , när det gäller budgetmässiga bestämmelser för centrala regeringar och regioner eller länder som är autonoma inom en stat ?
Jag skulle vilja svara MacCormick att kommissionen inte planerar att ändra bestämmelserna för additionalitet , som för perioden 2000-2006 anges i artikel 11 i den allmänna förordningen för fonderna .
Liksom i det förflutna anges det i dessa bestämmelser att additionalitetsprincipen skall tillämpas i förbindelsen mellan strukturfonderna och samtliga utgifter , jag säger utgifter , av medlemsstaten för utveckling .
I det avseendet måste man understryka att det är de utgifter som finansierats genom strukturfonderna som bör vara additionella .
Det krävs inte att samfinansieringen av medlemsstaten skall vara det , det vill säga läggs till de befintliga utgifterna .
Så länge som medlemsstaten inte minskar sina egna totala utgifter kan man anse och vi anser att strukturfonderna läggs till de nationella utgifterna och att additionalitetsprincipen således respekteras .
Vad beträffar de tillämpliga budgetbestämmelserna i medlemsstaterna mellan centralregeringen och regionerna eller i de länder som har en intern självständighet , bestäms de enbart utifrån nationella överväganden och berörs således inte av additionaliteten , i enlighet med förordningarna .
Jag ber om ursäkt för att ha gett detta ytterst juridiska svar .
Efter kontroll är det i varje fall på det sättet som vi rättsligt och exakt i förhållande till förordningen om strukturfonderna från Berlin bör definiera och förstå additionalitetsprincipen .
Jag är tacksam för ett tydligt svar men naturligtvis litet besviken på dess innehåll .
Vi har bara kvar artikel 11.1 som säger att anslag från fonderna får inte ersätta medlemsstaternas offentliga eller andra likvärdiga strukturella utgifter .
Nåväl : det skall vara den rådande regeln .
Tillåter artikel 11.1 möjligen följande praxis .
När en självstyrande region eller ett lands anslag från europeiska strukturfonderna ökar gör staten en åtföljande minskning av huvudfinansieringen till den regionen , så att det tillgängliga totala finansieringspaketet överensstämmer med en formel fastställd nationellt utan hänsyn till de strukturfondsmedel som beviljats av unionen .
Är det verkligen tillåtet ?
Tyvärr har jag inte tillräckligt med tid för att fördjupa mig och om herr MacCormick tillåter skulle jag vilja säga honom genom att ge honom delvis rätt i hans resonemang att jag kommer att komplettera mitt svar skriftligt och åter ge honom de rättsliga grunderna både för artikel 11 i allmänhet och artikel 11.1 i synnerhet .
Jag känner till , herr ledamot , med vilken kompetens ni följer alla dessa frågor .
Jag känner också till de särskilda problem som finns i ert valdistrikt i Skottland där vissa tvister eller diskussioner uppstår om dessa ämnen .
Jag påminner dock om att på ett allmänt plan är det utgifterna från strukturfonderna som skall vara additionella , enligt alla antaganden , och det är så att så länge som medlemsstaten inte minskar sina totala utgifter läggs strukturfonderna till de nationella utgifterna och vi anser att additionalitetsprincipen respekteras .
Jag skall ändå gå litet längre i mitt skriftliga svar som jag lovade er för att säga det mer objektivt och exakt .
Additionalitet är också en stor fråga i Wales , som jag företräder .
Senast förra veckan var den en av de frågor som förde fram till ett misstroendevotum mot och avgång av förstesekreteraren i nationalförsamlingen i Wales .
Så sent som 1991 och 1992 vann kommissionen en strid mot Förenade kungariket om additionalitet , vid tillfället kopplat till finansieringen från Rechar-programmet .
Detta ledde till att en överenskommelse undertecknades varmed Förenade kungarikets regering lovade att införa förfaranden för att se till att EU : s medel användes för de områden som de var avsedda och var i själva verket additionella medel .
Och ändå har vi fortfarande dessa problem i Wales och Skottland .
Kan kommissionen granska denna speciella situation mot bakgrund av den överenskommelse som undertecknades med Förenade kungarikets regering ?
Jag förstår således , fru ledamot , att den debatt som jag hade kännedom om i Skottland också pågår i Wales .
Jag skall kontrollera den punkt som ni anger och , om ni går med på det , kommer jag på samma gång att ge skriftligt svar på er fråga såsom jag lovade MacCormick .
Fråga nr 47 från ( H-0088 / 00 ) : Angående : Belopp som Andalusien kommer att få från strukturfonderna för perioden 2000-2006 Vilket belopp kommer Andalusien att få i bidrag från strukturfonderna för ovannämnda period enligt kommissionens uppskattningar och i enlighet med de kriterier som fastställdes vid toppmötet i Berlin , bland annat beträffande BNP per invånare , arbetslöshetsnivån och befolkningssiffran enligt 1996 års mantalslängd ?
Frågor till Bolkestein Jag skall anstränga mig , herr talman , att ge ett kort svar genom att säga till ledamoten att den regionala utvecklingsplan som lades fram av de spanska myndigheterna den 29 oktober gör det inte möjligt för mig att dra någon slutsats om en fördelning av gemenskapens medel mellan de spanska mål 1-områdena - eftersom det handlar om i Andalusien - och således de medel som var avsedda för den region som ni företräder .
Jag vill således säga er , fru ledamot , att eftersom jag inte lyckades se saken klart vände jag mig till ekonomi- och finansministern , Rato , med en skrivelse som jag har här från den 14 december för att be honom om vidare information om det framlagda dokumentet .
Under de kommande veckorna skall kommissionen inleda förhandlingar med de spanska myndigheterna för att utarbeta gemenskapsstödramen för den nya perioden 2000-2006 och vid dessa möten , det kan jag försäkra er , kommer kommissionen att få de nödvändiga klarläggandena om fördelningen per region .
Vad gäller Andalusien , kommer jag således att skynda mig att meddela er personligen , om ni vill det , så snart som jag förfogar över informationen per sektor och per region .
Herr kommissionär , problemet är att när Aznar vänder sig till Europeiska unionen för att ta betalt för samtliga andalusier , talar man om det för alla , men när Aznar skall betala i form av tjänster till den regionala regeringen i Andalusien , för samtliga andalusier , bortser han från fyrahundra tusen , och det är mycket allvarligt , för fyrahundra tusen barn är som om hela Strasbourg , eller en större stad som Granada , vore full av barn som Aznar inte ser .
Det är en viktig fråga och jag skulle vilja veta om herr kommissionär , för här kan man tala om barnbedrägeri , kommer att se till att andalusierna och Andalusien inte luras på dessa pengar , att de pengar som Europeiska unionen skall betala till Andalusien mot bakgrund av folkräkningen , inbegriper de fyrahundra tusen barn som Aznar inte räknar med när det gäller att förse dem med skolor och annan service .
Fru ledamot , jag vill be er alla - ta inte det här som en varning - att vi bara behandlar frågor som har med gemenskapen att göra .
Jag vet att dessa frågor är av stor betydelse i Spanien och det finns olika visioner ...
Jag kan påpeka för herr kommissionären att Aznar är Spaniens premiärminister .
Ni kan nu besvara frågan .
Fru ledamot , då jag hörde att ni har god röstkapacitet , hoppas jag att er röst var tillräckligt stark för att höras i Madrid , men jag förstod att det ni sade inte var riktat direkt till mig .
Jag har gett er mitt svar .
Jag är angelägen om att strukturfonderna , och särskilt de som rör mål 1 , skall delas ut där det finns behov .
Vi har kriterier som tillämpas och vi vet här indikativt vad varje område i Europa borde eller skulle kunna få .
Emellertid - jag gömmer mig inte bakom den , men jag är alltid tvungen att hänvisa till den allmänna förordningen , som jag bör diskutera med de nationella myndigheterna i varje land och med regeringen i varje land .
De har ansvaret att göra fördelningen så objektivt och rättvist som det är möjligt .
Jag behöver veta i alla fall och därför sade jag att jag inte kan svara i dag .
Eftersom jag inte har svaret , skrev jag till ekonomi- och finansministern den 14 december .
Nu kommer den tid då jag blir otålig över att inte ha fått svar , men jag kommer att vidarebefordra det till er när jag får det .
Jag beklagar att herr kommissionären än en gång har blivit delaktig i en fantasirik och i det här fallet lidelsefull inblandning .
I Spanien - det vill jag påminna er alla om - befinner vi oss inte bara i valtider , det är tjugofem dagar kvar till valet .
Det är en tröst för kommissionären att valen kommer att äga rum om tjugofem dagar , för sedan är det troligtvis ingen som kommer att ställa den här typen av frågor till honom längre .
Jag tycker verkligen att det är viktigt att tala om att Andalusien kommer att få 50 procent mer inom gemenskapens ramar och att Spanien dessutom slår rekord vad gäller att förverkliga strukturfonderna , något som innebär att fördelningen sker helt i enlighet med tillämpningsbestämmelserna , att den är decentraliserad och att den ske enligt planerna för regional utveckling och de olika ramarna för gemenskapsstöd .
Som en avslutning vill jag ställa en konkret fråga till herr kommissionären : Anser ni att tillämpningsbestämmelserna för strukturfonderna bör ändras eller anser ni att de nuvarande fördelningskriterierna är godtagbara ?
Jag tycker att debatten är mycket spännande .
Jag förstår väl att den har en dimension som inte endast gäller gemenskapen .
Därmed sagt att vi måste tänka på att det ständigt är val i samtliga unionens länder .
Det som är mig ett nöje det är att strukturfonderna i grunden är ett diskussionsämne i Grekland och i Spanien .
Nyss talade vi här om medborgardebatt och offentliga debatter .
Desto mer man talar om Europa och det som Europa gör för det dagliga livet , även om man grälar litet , ju bättre är det , förutsatt att man talar om det objektivt .
Jag skall inte säga vad jag känner , herr ledamot , om en eventuell förändring av förordningen om strukturfonderna .
Den antogs just i Berlin i förra året .
Jag genomför den för de kommande sex åren .
Vi kommer att tala om den med anledning av betänkandet om sammanhållning som är ett viktigt möte för mig här , med er , och inför er , för att göra en sammanfattning och på samma gång dra upp riktlinjer , och det ögonblick kommer i början av nästa år , då vi skall ta upp eventuella justeringar och eventuella ändringar .
Jag ber er , låt mig just nu tillämpa den förordning som ännu inte tillämpats , eftersom den är daterad i Berlin .
Det är vad jag kan säga i dag .
Tack så mycket , herr Barnier , för era svar .
Frågorna 48 till 50 kommer att besvaras skriftligen .
Fråga nr 51 från ( H-0049 / 00 ) : Angående : Nya lokaler för Byrån för harmonisering inom den inre marknaden För närvarande fortsätter Byrån för harmonisering inom den inre marknaden att arbeta i sina gamla provisoriska lokaler trots att den nya byggnaden invigdes i juni 1999 .
Dessa ovanliga omständigheter motiverar följande fråga till kommissionen : Vilka är orsakerna till att Byrån för harmonisering inom den inre marknaden ännu inte flyttat in i de nya lokalerna ?
Ledamoten ställde en fråga i det här ämnet i november 1999 och jag skulle gärna vilja hänvisa till det svaret .
Dessutom har jag med anledning av den nya frågan bett ordföranden för Byrån för harmonisering inom den inre marknaden , Alicante-byrån alltså , om en kommentar och jag kan därför för byråns räkning meddela ledamoten följande : Byrån är ännu inte klar att flytta in i den nya byggnaden .
Tyvärr har vissa tidsfrister överskridits .
Ett antal tekniska arbeten återstår , till exempel ett datornät , arkivutrymmen , en restaurang och möbler .
Harmoniseringsbyrån håller på med detta och räknar med att flyttningen till den nya byggnaden skall kunna ske i juni .
Föregående fråga föranledde oss att tala om valen .
Jag tror att saken kom upp i samband med den frågan för ni , herr kommissionär , var inte med på den så illusoriskt kallade " officiella invigningen " av sätet för Byrån för harmonisering inom den inre marknaden den 9 juni , mitt under valkampanjen , och sådana äger inte bara rum i Spanien inför Europavalen utan även inför de lokala och regionala valen .
Om ni hade varit där , skulle ni garanterat ha tyckt att det var pinsamt .
Kommissionens ordförande och några kanslichefer var visserligen på plats .
Mitt under pågående valkampanj höll flera auktoriteter , alla från regeringspartiet , några anföranden som var uppenbart valfläsk och som dessutom direktsändes i TV .
Synnerligen märkligt var anförandet av Valencias regionalpresident som ägnade sig åt att lovorda den spanska regeringens liksom den egna regionala regeringens insatser , något som inte alls hörde till saken .
Att mitt under pågående valkampanj inviga en byggnad som inte är färdig , och som åtta månader efter invigningen inte har kunnat användas , har skapat en ytterst pinsam situation för den spanska regeringen .
Det bekymrar mig inte att den spanska regeringen har gjort bort sig , för när allt kommer omkring är det deras ansvar , däremot bekymrar det mig att kommissionen gör det genom att med sin närvaro garantera ett sådant icke representativt agerande .
Därför vill jag fråga er , herr kommissionär : Finner ni det normalt att inviga en byggnad mitt under en valkampanj innan den ens är färdig ?
Finner ni det normalt att kommissionen genom sin närvaro garanterar ett sådant icke representativt agerande från den spanska regeringens sida ?
Det hör inte till mina uppgifter att uttala mig om inrikespolitiska situationer i den ena eller den andra medlemsstaten .
Därför vill jag heller inte kommentera den situation som Berenguer nyss tog upp .
Jag måste erkänna att jag inte känner till av vilken anledning en viss öppningshögtid i Spanien äger rum .
Jag kan dock säga att jag hoppas att den här byggnaden äntligen skall tas i bruk så snart som möjligt .
Vidare vill jag tala om att jag själv hoppas att vara närvarande i Alicante i slutet av maj för att tala vid en konferens där .
Jag hoppas att byggnaden då skall ha tagits i bruk .
Jag vill påpeka för kommissionären att det inte rör sig om en valfråga .
Som medlemmar av utskottet för rättsliga frågor och den inre marknaden har vi sett hur denna institution har skapats och det är uppenbart att den invigdes av valmässiga skäl .
I dag - ett år senare - har den fortfarande inte tagits i bruk , och det innebär att kommissionen använde pengar på en falsk invigning .
Man kan gott fråga sig om en användning av medel till en falsk invigning var motiverad .
Ännu en gång , kommissionen håller sig inte sysselsatt med skälen till olika handlingar i medlemsstaterna .
Kommissionen bryr sig om det som tillkännages offentligt och vad som görs .
Vi tänker inte ge oss in i något som på franska kallas un procès d ' intention .
Vi bryr oss om offentliga , officiella handlingar och händelser och inte eventuella bakomliggande motiv .
Därför tycker jag också att det i det här fallet är svårt att svara Medina på hans fråga .
Kommissionen undrar inte över av vilken anledning något sker tidigare eller senare , förutom att kommissionen uppskattar att en byggnad , som för den här byrån , öppnas och tas i bruk så snabbt som möjligt .
Vidare håller sig kommissionen inte heller sysselsatt med om vissa utgifter skedde reellt eller virtuellt .
För min del är alla utgifter reella .
Vidare låter jag historien vara som den är .
Eftersom frågeställaren är frånvarande , bortfaller fråga nr 52 .
Eftersom de behandlar samma ämne , kommer frågorna 53 och 54 att tas upp tillsammans .
Fråga nr 53 från ( H-0057 / 00 ) : Angående : Svenska undantagsregler vad gäller införsel av alkoholhaltiga drycker över gränsen Sverige har i dag ett undantag till år 2004 som medger en begränsning av alkoholhaltiga drycker över gränsen .
Svenska regeringen och en stor folkopinion har uttryckt att detta undantag måste förlängas av folkhälsoskäl .
Kan kommissionen redogöra för sin inställning till det svenska undantaget beträffande införsel av alkoholhaltiga drycker ?
Fråga nr 54 från ( H-0117 / 00 ) : Angående : Alkoholmonopol och den inre marknaden Vilka åtgärder avser kommissionen att vidta för att förhindra den förlängning av det statliga alkoholmonopolet som Sverige uppenbarligen planerar , och de införselrestriktioner som följer därav , samt för att se till att den inre marknadens bestämmelser får genomslag ?
Jag skulle vilja besvara de här två frågorna på följande sätt .
Vid tillträdet till Europeiska unionen fick Sverige behålla de kvantitativa begränsningarna för alkoholhaltiga drycker som resenärer får föra in i landet från andra medlemsstater .
Det här undantaget från principen om fri rörlighet för varor och personer slutar att gälla den 30 juni i år .
Sverige vill nu ha en förlängning av den här åtgärden i ytterligare fem år eftersom det skulle vara nödvändigt för att skydda folkhälsan .
Min inställning i den här frågan är tydlig .
Sverige har nu haft tillräckligt god tid på sig sedan anslutningen till unionen för att anpassa sin politik till ett tillstånd utan sådana importrestriktioner .
Därför ser jag inget skäl till varför jag skulle föreslå en förlängning av det här undantaget .
Europeiska medborgare har rätt att för egen räkning köpa varor inklusive skatter , i vilken medlemsstat de vill och sedan ta med dessa varor till en annan medlemsstat utan att de här varorna måste genomgå kontroller och utan att nya skatter eventuellt måste betalas .
Det är en grundprincip för den inre marknaden och avvikelser från den principen måste vara undantag och tidsbegränsade .
Vi vill garantera att svenska medborgare nu också skall kunna åtnjuta fördelarna med den inre marknaden , precis som andra medborgare i Europeiska unionen kan göra .
Det betyder inte alls att jag inte delar oron i Sverige angående de möjliga hälsoproblem som kan förorsakas av alkoholmissbruk .
En undersökning som nyligen gjordes av professor Lindgren vid universitetet i Lund visade dock att ett avskaffande av begränsningarna inte skulle leda till en högre alkoholkonsumtion i Sverige .
Jag har redan vid två tillfällen kunnat diskutera min hållning med Bosse Ringholm , Sveriges finansminister .
Förra veckan diskuterade jag också den här frågan med den svenska riksdagens finansutskott .
Det är nu upp till den svenska regeringen att vidta lämpliga åtgärder .
Tack för svaret , herr kommissionär .
Jag vill bara beklaga att det står fel i min fråga till kommissionen .
Det står nämligen år 2004 , men det skall naturligtvis vara den 1 juli år 2000 .
Jag har till viss del förståelse för kommissionens ståndpunkt att undantag skall vara tillfälliga .
Det är en regel som är normal .
Ändå skulle jag vilja ställa två frågor : Tänker ni ändå ta upp fortsatta diskussioner med den svenska regeringen om en förlängning av undantagen , exempelvis så länge som Danmark och Finland har undantag ?
Min andra fråga handlar om den samlade alkoholpolitiken .
Man kan ju se detta som en fråga rörande den inre marknaden , men också som en folkhälsofråga för hela EU .
Vilken roll spelar alkoholpolitiken i kommissionens arbete , och vilken roll spelar folkhälsoaspekterna ?
Alkoholpolitiken i hela Europa handlar inte bara om den inre marknaden , utan också om folkhälsan .
Hade vi totalt sett betraktat dessa aspekter , hade det kanske varit lättare att föra diskussionen med Sverige .
Får jag be att få tacka herr Andersson för fortsättningen på hans första fråga och den frågan vill jag svara på så här .
För det första så har Finland och Danmark undantag från grundregeln om fri rörlighet för varor fram till år 2003 .
De länderna håller på att vidta förberedande åtgärder så att de är klara för fri tillgång till alkoholhaltiga produkter år 2003 .
När det gäller Sverige så är situationen litet annorlunda .
Där beslutade man 1995 om en undantagsperiod på fem år och den går ut nu .
Jag har ännu inte hört några argument som skulle kunna ligga till grund för att kommissionen borde förlänga den perioden .
För det andra så förs ständiga förhandlingar med den svenska regeringen .
Jag kan meddela Andersson att jag måndagen den 6 mars reser till Stockholm för att där samtala med minister Ringholm , med svenska riksdagsledamöter och om så önskas även med statsministern eller med andra ministrar , för att prata vidare om den här frågan som - det inser jag helt och fullt - ger anledning till starka politiska känslor i Sverige .
För det tredje så förstår jag naturligtvis mycket väl att hälsoaspekten av den här frågan är viktig .
Jag upprepar för andra gången att professor Lindgren vid universitetet i Lund har sagt att , vad som än sker med avseende på importbegränsningarna , alkoholkonsumtionen i Sverige kommer att ligga kvar på samma nivå .
Frågan är då naturligtvis var den mängd alkohol som inte förs in av resenärer då kommer ifrån .
Svaret är att den antingen smugglas in eller också tillverkas den av svenska invånare själva och som Andersson vet så är det ett mycket farligt och ohälsosamt förfarande .
Andersson verkar tro att hälsosituationen går framåt om vi begränsar importen av alkohol .
I det fallet skulle inte bara Sverige , utan alla länder i Europeiska unionen vara tvungna att utgå från principen att all försäljning av alkohol skall förbjudas .
Vi hade ett sådant exempel i Förenta staterna .
Andersson känner säkerligen till det som då kallades för prohibition .
Han vet också vilka följder det hade för maffians verksamhet i Förenta staterna , där man slutligen också gjorde slut på denna prohibition .
Allt det här betyder att man naturligtvis måste skydda hälsan men inte genom att förbjuda alkohol , det hjälper nämligen inte .
Herr talman !
Det handlar ju i verkligheten om intäkter från det svenska alkoholmonopolet , och om den svenska regeringen säger att den måste använda dem för att täcka kostnader för hälsovården , så är detta ändå ett bevis för att det innebär en snedvridning av konkurrensen , ty andra länder måste själva finansiera sina hälsovårdskostnader , utan att förfoga över något alkoholmonopol .
Min fråga gäller om ni också känner till undersökningar om att en måttlig konsumtion av alkohol av hög kvalitet , alltså exempelvis frankiskt vin eller bayerskt öl , rent av är hälsofrämjande , och att det därigenom rent av skulle ske en avlastning av den svenska statsbudgeten ?
Om jag förstått det rätt så har Posselt börjat peka på skatteaspekterna av den här frågan .
Jag tror mig också veta att den höga skatten på alkoholhaltiga drycker i Sverige har sitt ursprung år 1638 och att staten sedan dess får en ansenlig del av sina skatteinkomster från försäljningen av alkoholhaltiga produkter .
Som ni vet så är det nu ett statligt monopol i Sverige , vilket i sig inte heller är helt i enlighet med EU-lagstiftningen .
När det gäller alkoholens hälsosamma verkan - för jag tror att Posselt talade om det också - så är jag helt ense med honom : jag tror att en bra flaska vin kan vara mycket bra för hälsan och socialt sett dessutom mycket angenäm .
Kanske kan Posselt , Andersson och jag själv träffas i parlamentets bar en dag och dricka en akvavit tillsammans .
Herr talman !
Jag lyssnade med intresse till kommissionärens svar på kravet att tillämpa den inre marknadens bestämmelser .
Jag undrar om han kan säga om han anser sitt svar vara i överensstämmelse med kommissionens underlåtenhet att dra den franska regeringen inför EG-domstolen avseende tillämpningen av Frankrikes " Loi et Vin " , som effektivt hindrar den inre marknadens bestämmelser att gälla vid försäljning av alkohol och alkoholprodukter i Frankrike ?
Kan vi nu förvänta oss att Europeiska kommissionen vidtar åtgärder mot den franska republiken hos EG-domstolen ?
Jag skulle vilja kort besvara den fråga som ställdes av ärade ledamoten eftersom detta ärende nu är under övervägande hos kommissionen .
Kommissionen måste fatta ett beslut om ärendet är avslutat eller om det skall hänskjuta det till EG-domstolen .
Mitt svar är kanske inte tillfredsställande just nu , men jag lovar den ärade ledamoten att kommissionen skall fatta det beslutet inom några veckor .
Jag ber om ledamöternas förståelse för denna lilla försening av kommissionens beslut .
Herr kommissionär !
Har ni något skäl med hänsyn till folkhälsa till en skillnad i skattesats för till exempel , skotsk whisky eller franskt bordeauxvin eller mina kollegors bayerska öl ?
Kan ni tänka er en likvärdig grund alkoholbeskattning i Europa ?
Frågan om punktskatter som den ärade ledamoten hänvisar till är den berörda medlemsstatens prerogativ .
Kommissionen har inga medel att genomdriva någon särskild minskning eller ökning av punktskatter på alkoholprodukter eller några andra produkter .
Mot slutet av detta år kommer kommissionen att överlämna en rapport om skillnaderna i punktskatter mellan medlemsstater .
Den kommer utan tvivel att leda till diskussioner både med parlamentet och rådet om det nuvarande läget i denna fråga , vilket tyder på att det finns ganska stora skillnader i punktskattesatser mellan medlemsstater .
Exempelvis , och jag tror att den ärade hänvisade till detta , tillämpas inga punktskatter på vin i Frankrike medan de tillämpas i Förenade kungariket .
Det leder till en snedvridning av den inre marknaden eftersom vin smugglas från Frankrike till Förenade kungariket .
Frågan gäller i synnerhet förhållandet mellan punktskatter och alkoholhalten i de varor som är punktskattepliktiga .
Kommissionen har inga möjligheter att påverka i denna fråga .
I Sverige används punktskatter rent av för att minska alkoholkonsumtionen .
Även om detta leder till en skillnad i punktskattesats mellan Sverige och andra medlemsstater i unionen - och det i sig självt ökar gränssmugglingen av alkoholprodukter - är det ett lagligt instrument för att minska alkoholkonsumtionen .
Det finns naturligtvis efterfråge-elasticitet , i detta fall efterfråge-elasticitet rörande pris .
Jag är inte exakt säker på vad det är men det är inte noll , därför bör den ge någon effekt .
Min fråga skulle ha blivit nästan exakt den som Purvis ställde , men jag skulle vilja gå vidare i frågan .
Förutsatt , som ni säger , att punktskatter är medlemsstaternas prerogativ , kan ändå användning av det prerogativet på ett sätt som är diskriminerande mot producenter i en del av gemenskapen till skillnad mot andra fortfarande strida mot den inre marknadens princip .
Om vi till exempel tar vad Purvis och jag skulle tänka på , de maltwhiskyproducerande delarna av skotska högländerna - ett verkligt ytterområde i Europa med hårda ekonomiska villkor , ett helt lantbrukssamhälle liksom ett destilleringssamhälle beroende av detta - en generell praxis att beskatta alkoholen i skotsk whisky , holländsk gin eller dansk akvavit mer än alkohol i öl eller vin tycker jag verkar diskriminerande och en diskriminerande tillämpning av något som onekligen ligger inom medlemsstaternas prerogativ .
Får jag försäkra MacCormick och övriga ledamöter av detta parlamentet att den nuvarande situationen med punktskatter som skiljer sig mellan medlemsstater är verkligen något som inte är bra för den inre marknadens funktion .
Vi måste begränsa oss till alkoholprodukter .
Om man ser på olja till exempel finner man att punktskattesatserna i Tyskland skiljer sig från dem i Holland och följaktligen åker holländska motorister över gränsen och tankar i Tyskland .
Det är i själva verket en snedvridning av den inre marknaden .
Om jag fick göra som jag ville skulle jag svänga en trollstav och likställa alla punktskatter i hela Europa .
Följden skulle bli att smuggling upphörde utom i de fall produkter var väsentligt dyrare i en medlemsstat än i en annan .
Men jag har inget trollspö och jag får inte göra som jag vill .
Detta är ett område för enhällighet , som MacCormick vet , och om inte alla medlemsstater går med på att likställa punktskatter , kommer det inte att ske .
Ännu en gång , mot slutet av detta år kommer kommissionen att överlämna en rapport om det nuvarande läget rörande punktskatter och jag finns naturligtvis tillgänglig för diskussioner med parlamentet om den rapporten .
Tack så mycket herr kommissionär .
I dag kommer vi att följa ert råd och dricka ett - eller kanske två - glas vin från Alsace .
Vi vet inte vilka pålagor det vinet har , men jag förmodar att även det är belagt med höga skatter .
Eftersom tiden för frågor till kommissionen är ute , kommer frågorna nr 55 till 114 att besvaras skriftligen .
Jag förklarar härmed frågestunden med frågor till kommissionen avslutad .
( Sammanträdet avbröts kl .
19.30 och återupptogs kl .
21.00 )
 
Gemenskapsåtgärder på vattenpolitikens område ( fortsättning på debatten ) Nästa punkt på föredragningslistan är fortsatt debatt om andrabehandlingsrekommendationen om gemenskapsåtgärder på vattenpolitikens område .
Herr talman !
Situationen för Europas sötvatten är inte lika allvarlig som i andra del av världen , men rent allmänt är det ett bevisat faktum att efterfrågan på vatten ständigt ökar samtidigt som kvaliteten minskar .
Därtill kommer de problem med förorening av vattnet som de potentiella nya medlemsstaterna i öst tampas med .
För övrigt har en behållare med cyanid just gått sönder i Rumänien , något som utgör ett hot mot grundvattenakviferer som förser Jugoslaviens befolkning med vatten .
Jag har förstått det som att Wallström , vars närvaro här i kväll jag uppskattar , kommer att besöka området .
Jag tror inte att något land , någon regering och givetvis inte någon medlem av parlamentet kan låta bli att erkänna behovet av detta direktiv för att sätta stopp för den nuvarande uppdelningen av vattenpolitiken och underlätta igångsättandet av ett program med specifika åtgärder för olika vattendrag .
Det har varit svårt och komplicerat att ta fram direktivet , det är många intressen som står på spel och åsikterna är delade .
Jag tvivlar inte på att den här mandatperiodens föredragande , Lienemann , har lagt ned stor möda och stort engagemang på att förena och återförena olika ståndpunkter , och hon har i stor utsträckning lyckats med det .
Däremot är det nästan omöjligt att känna till och rättvist bedöma alla situationer och förväntningar .
Jag kommer från ett land vars södra del vetter mot Medelhavet och där tillgången till vatten historiskt sett har berott på växlingarna i ett ombytligt klimat och markens svåra beskaffenhet .
I Medelhavsområdet har man varit tvungen att kämpa för sin utveckling genom att sträva efter att övervinna dessa svårigheter sekel efter sekel , år efter år , dag efter dag fram tills i dag .
Som viktig betraktar vi därför direktivets praktiska tillämpning av den skyldighet som fastslås i artikel 164 i fördraget angående att i gemenskapslagstiftningen skall hänsyn tas till regionernas mångfald .
I tillämpningen av just denna princip protesterar den spanska delegationen i Europeiska folkpartiet mot ändringsförslagen 4 - stycke 21 - , 13 och 49 - artikel 11d ) - , eftersom de utgör starka begränsningar på ett område som är medlemsstaternas , nämligen regleringen av vattenresurserna .
Det skulle vara mycket svårt för gemenskapen att fastställa villkoren för reglerandet av dessa i de olika regionerna , med tanke på den interna balans som alltid står på spel och som under alla omständigheter kräver goda kunskaper om de olika områden och intressen som berörs .
Likaså förkastar vi de ändringsförslag enligt vilka man vill inbegripa den totala vattenkostnaden år 2010 .
Det råder ingen tvekan om att vi måste fastställa vattenpriser som främjar en effektiv användning , men som samtidigt gör att konkurrenskraften bevaras inom de produktiva sektorerna i de minst gynnade regionerna och inte hindrar en rättmätig utveckling .
Slutligen vill jag nämna något angående ändringsförslagen om farliga ämnen , där det fastslås att en nollgradig eller nära nollgradig förgiftning skall uppnås .
Hittills har ingen nollgradig förgiftning upptäckts i samband med mänskliga aktiviteter .
Mina damer och herrar , vi kommer inte att göra målen i detta viktiga direktiv rättvisa om vi inte kan förse det med den flexibilitet och anpassbarhet som krävs för att garantera att direktivet uppfylls .
Jag hoppas att parlamentet än en gång röstar utifrån verkligheten och med respekt för subsidiaritetsprincipen och söker uppnå en bra jämvikt mellan miljömålen och de ekonomiska och sociala hänsynen , de tre viktiga komponenterna för att uppnå en hållbar utveckling som vi alla så gärna vill ha .
Herr talman , ärade kommissionär !
Detta är ett mycket viktigt direktiv .
Målsättningen är ju att förbättra vattenkvaliteten och säkerheten i vattenförsörjningen .
Medborgarna måste ha rätt till rent vatten .
Det är viktigt för såväl miljön som för folkhälsan .
Jag talar inte alls för egen del , eftersom jag händelsevis råkar höra till de få lyckligt lottade européer som kan dricka vatten direkt från den egna sjön .
Vi måste se till att vi snabbt kommer igång med att förbättra vattenkvaliteten .
Vi måste genast börja arbeta på det .
Vi har inte råd att vänta .
Det är viktigt att tidtabellen är ambitiös .
Jag anser det inte vara för ambitiöst om vi utgår ifrån att vi år 2020 inte längre släpper ut föroreningar i vattnen och att vi strävar efter att till dess uppnå en nollnivå när det gäller föroreningar och giftiga ämnen .
Det är ju fråga om att vi gör det som är tekniskt möjligt ; mer än så kan det ju inte vara frågan om , men vi måste vara tillräckligt ambitiösa .
Jag vill göra er uppmärksamma på en sak som också har diskuterats tidigare .
Jag anser att utskottet för miljö , folkhälsa och konsumentfrågor alltför snävt avgränsat frågan om transport av vatten .
Detta är inte enbart Spaniens problem , det är också de nordiska ländernas problem och jag hoppas verkligen att man i dessa frågor förlitar sig på nationella lösningar då dessa miljömässigt och ekonomiskt sett är bättre än de som nu framförs i direktivet .
Herr talman , fru kommissionär !
Grattis , Lienemann , till ett utmärkt arbete !
Vatten och luft omger oss överallt .
Vi delar dem med alla människor på denna jord .
Vatten är en förutsättning för mänskligt liv .
Och vi blir alltfler som lever i detta liv .
Schleicher antydde tidigare i dag att det skulle vara orealistiskt med rent vatten .
Ingenting kan vara mer fel !
Det är orealistiskt att successivt försämra vattenkvaliteten , att successivt försämra livsförutsättningarna .
Särskilt orealistiskt är det för jordbruket , som är mest beroende av en ren natur och rena resurser .
Därför vill jag vädja till parlamentets ledamöter att inse att hårda krav på en ren miljö innebär den största realismen på lång sikt .
Herr talman !
Både vi och jag personligen stöder Leinemanns betänkande , de mål det uppställer och det direktiv vi diskuterar .
Vi borde emellertid försöka se litet längre .
T.ex. i mitt land , herr talman , är det ett gigantiskt problem att man ändrar flodernas lopp och torrlägger sjöar med stöd av ihåliga argument och naturligtvis med stora risker både för grundvattnet och för ytvattnet .
Även om vi kommer fram till vem som beslutar om sådana ingrepp , anser jag att vi behöver gemensamma och mycket stränga regler .
Det stora problemet , fru kommissionär , är dock enligt min mening planeringen för att återställa grundvattenreserverna och flodernas naturliga lopp och att åter fylla sjöarna med vatten .
Detta måste ske under de tio år som vi planerar för .
Jag anser att man måste kunna välja och finansiera sådana projekt , eftersom de kan ha en utomordentligt stor betydelse för utvecklingspolitiken .
Herr talman !
Här har vi något som i grunden är ett bra åtgärd .
Den lägger fast uppnåbara normer grundade på subsidiaritetsprinciper och förvaltning av vattenresurser .
Dess syfte med bra dricksvattenkvalitet , för djur- och växtliv , miljön och för ekonomiska ändamål är rätt .
Att förhindra miljöförstöring och vattenförsämring måste vara rätt liksom möjlighet att förvalta vattenresurser vid torka och översvämning .
Vi har tre olösta problem .
Det första är ledning av vatten mellan vattenområden .
Det är en fråga som berör mina kollegor från Spanien , Irland och Förenade kungariket .
Ändringsförslagen 4 , 49 och 87 kan inte godkännas eftersom de skulle begränsa möjligheten för ett land att leda vatten från där det finns till där det behövs , vare sig det gäller områden med torka eller städer .
För det andra måste vi ha realistiska mål , men målsättning i alla fall .
Om man granskar ändringsförslag 7 till exempel , som kräver fullständigt avlägsnande av naturligt förekommande ämnen , kan ni inse att några av de uppställda målen är orealistiska .
Vidare är några av målen satta till nästan noll - på engelska är det en ganska meningslös term .
Vi måste granska dessa mycket noga .
Konceptet att fortsätta minskningen , såsom i ändringsförslag 58 , är mycket bättre .
För det tredje tar jag upp problemet för skotsk whisky .
Skotsk whisky - särskilt maltwhisky , som är den bästa - kräver vattenextraktion som används till en viss mängd och sedan återförs till vattensystemen .
En del av det slutar i flaskan och dricks upp .
Vi måste se till att man i ändringsförslag 49 och 87 tar bort undantaget om att den skall utgå så att whisky kan fortsätta att drickas som " high quality " , vilket innebär att man för den måste använda bra , skotskt torvvatten .
Det är min tredje begäran - att vi granskar noggrant dessa åtgärder innan man godkänner hela denna åtgärd .
Herr talman , ärade kollegor , fru kommissionär !
Det ramdirektiv vi i dag granskar i en andra behandling är en slags grundlagsenlig skrivelse som berör allt från vatten till Europeiska unionen .
Direktivet utgör på en och samma gång såväl ankomst som avresa .
Ankomst därför att det förbereddes av ett helt batteri av direktiv , dock fragmentariska och utspridda , som lämnade spår av logisk helhet och systematiskt sammanhang när det gäller lagstiftning om vatten .
Det är också en avresa eftersom nya referensramar skapas som den framtida europeiska lagstiftningen om vatten skall anknyta och härledas till .
Ramdirektivet utger sig för att vara ambitiöst och realistiskt , voluntaristiskt och genomtänkt , vilket mer än väl uppnås .
De ändringsförslag som lades fram av kommissionen , tack vare ledamot Lienemanns utmärkta arbete , är till för att förstärka texten i direktivet och göra den mera rigorös .
Att göra den mera rigorös betyder inte att den blir mindre flexibel , om man bortser från de klimatologiska och geografiska skillnader som är så flagranta på europeiskt territorium .
Jag stöder till fullo förslaget till betänkande , så tillåt mig applådera det samtidigt som jag vill säga att det finns två saker som oroar mig .
Först och främst en applåd : Enligt min mening är det ett oförnekligt framsteg att man i direktivet ställer krav på en integrerad förvaltning av hydrografiska flodområden och att vattenöverföringen mellan dessa områden bara skall göras när det visar sig vara absolut nödvändigt .
På till exempel Iberiska halvön är detta en hälsosam och pedagogisk princip till exempel på Iberiska halvön. är enligt min mening Min första oro gäller direktivets tidsplan : Den kan visa sig bli svår att följa , även om jag också tycker att det är en stor utmaning .
Min andra oro kan ni kanske gissa er till : Det kommer att bli svårt att fastställa kostnaderna för vattnet och bestämma respektive pris , särskilt när miljökostnaderna tillkommer , något som främst bland jordbrukarna framkallar misstro .
Att betala ett rättvist pris för vattnet kan också generera orättvisor .
Ramdirektivet är i sig en stor vadhållning : att europeiskt vatten år 2020 skall vara återställt till sitt ursprungliga skick , fri från föroreningar och utan farliga substanser .
En utopi ?
En återgång till det förindustriella samhället ?
Jag tror inte det .
Jag har fullt förtroende och känner stor optimism för det här .
Den katastrof som nyligen inträffade vid Donau kan , som i en mardröm , illustrera att en långsiktig politik och strategi för ett ekologiskt skydd av vattenområdena , oavsett vad det kan kosta , inte är de rikas lyx utan civilisationens absoluta nödvändighet .
Herr talman !
Först vill jag påtala det bottenlösa hyckleriet hos dem som , samtidigt som de skryter om sitt engagemang för miljön och för vattnet , gör sig skyldiga till så brottsliga handlingar som attackerna mot Jugoslavien , attacker som inte bara resulterat i tusentals döda och sårade utan också lett till ekologiska katastrofer när det gäller vattenreserverna , genom att vattnet inte bara blivit obrukbart utan också utomordentligt skadligt .
I anslutning till betänkandet skulle jag också vilja säga att principen om kostnadstäckning för vattenmyndigheterna absolut inte får tillämpas så att den leder till ökad beskattning av de ekonomiskt svagaste befolkningsgrupperna eller till att de små och medelstora jordbruken slås ut på grund av de enorma kostnaderna för bevattning .
Jag vill också påpeka att speciellt i områden med akut vattenbrist som i mitt land , i synnerhet på öarna , är det absolut nödvändigt att ge bidrag till investeringar i infrastruktur .
Syftet är att man skall spara på vatten , inte genom prisökning utan genom att öka tillgången på vatten framför allt genom att ta till vara det regnvatten som i dag rinner bort till ingen nytta och på sin väg till havet eroderar marken med alla de problem som detta innebär .
Därför stöder jag ändringsförslag 107 av vår kollega Marset Campos .
Dessutom är det nödvändigt att ta till vara flodvattnet bättre för att garantera fortsatt liv i områden som ständigt lider brist på vatten .
Slutligen vill jag säga att det är omoraliskt av rådet att , i likhet med kommissionen , påstå att det inte behövs många konkreta hänvisningar och förtydliganden , eftersom de täcks av exemplen i direktivet eller behandlas i andra delar av direktivet .
Syftet är att man vill behålla ett till hälften insynsskyddat område , vilket innebär att man under den första perioden , då direktivet tillämpas slutgiltigt , kan fatta en hel del avgörande beslut till gagn för storkapitalet .
Herr talman !
Jag vill först och främst säga att just skyddet av vattenmiljön , både vad gäller yt- och grundvattnet , förmodligen är ett av våra allra viktigaste åtaganden .
Det är det för att vi kan säkerställa tillräckliga vattenresurser , men också i hög grad för att skydda vattenresurserna mot föroreningar , så att vi även i framtiden skall få rent dricksvatten .
Att ha tillgång till rent dricksvatten är en rättighet för oss alla .
Jag vill gärna uttrycka ett stort erkännande av Lienemanns arbete i denna fråga .
Hon har utfört ett kolossalt arbete och jag vill gärna ge mitt stöd till alla Lienemanns ändringsförslag , som alla förbättrar den gemensamma ståndpunkten .
Och jag skall bara betona det viktigaste .
Först och främst tycker jag det är viktigt att vi fastställer vissa tydliga målsättningar för vattnets tillstånd redan före en period på tio år .
Jag tycker också att det är viktigt att vi utövar påtryckningar på medlemsstaterna så att de utarbetar de nödvändiga åtgärdsprogrammen snabbare än vad som uttrycks i den gemensamma ståndpunkten .
Slutligen vill jag säga att jag tycker att de åtstramningar som sker med hänsyn till betalningssystemen och prisfastställandet är korrekta , så att vi som konsumenter snabbare får en effektiv användning av vattenresurserna och samtidigt ett system som kan främja uppfyllandet av de miljömål som jag tror det råder stor enighet om .
Även här tycker jag att tidsfristen fram till år 2010 är en lämplig tidsfrist .
Slutligen vill jag säga att jag tycker det är mycket viktigt att vi kan inleda den gradvisa reduceringen av utsläpp av farliga ämnen .
Att vi kan göra det gradvist , men att vi samtidigt fastställer ett slutligt mål , dvs. år 2020 , när vi förhoppningsvis är nere på obefintliga utsläppsnivåer .
Om det inte är möjligt att fastställa detta som mål , är jag naturligtvis beredd att stödja det förslag som avser att vi skall nå mycket nära noll under år 2020 .
Jag tycker att Lienemanns förslag utgör en bra grund för vidare förhandlingar med rådet .
Herr talman !
Jag vill tacka föredraganden av betänkandet för ett förtjänstfullt arbete i beredningen av ett viktigt direktiv .
Den andra behandlingen av vattendirektivet kommer vid en läglig tidpunkt : De skakande nyheterna från miljökatastrofen i Rumänien måste utnyttjas både i dagens debatt och då man mera allmänt dryftar miljödimensionen i samband med utvidgningen av unionen .
Allra först måste man hitta de skyldiga till dådet och ställa dem till svars .
Cyaniden och tungmetallerna som hamnat i floden är fruktansvärda exempel på hur en vårdslös inställning till miljön kan fördärva vattendragen i tiotals år framöver .
Händelsen visar att miljönormerna och inställningen till miljön i några av de länder som ansökt om EU-medlemskap ännu befinner sig ljusår från EU-nivån .
Det vore också bra om unionen än en gång övervägde hur stöden till miljöprojekt skulle kunna styras för att stödja en hållbar vattenpolitik .
Med tanke på förslaget till direktiv är det bekymmersamt att man under granskningarna i utskottet för miljö , folkhälsa och konsumentfrågor inte tillräckligt beaktar de oförorenade ytvattnens betydelse för de naturliga grundvattenförekomsternas utbredning .
I Finland är ytvattnen mycket rena .
Tillverkningen av så kallat konstgjort grundvatten är ett ekologiskt sätt att filtrera rent ytvatten som påfyllning till grundvattenreserverna .
Processen kräver inga kemiska reningsverk .
Direktivet får inte äventyra denna verksamhet .
Utskottet för miljö , folkhälsa och konsumentfrågor försöker också genom att avvika från rådets gemensamma ståndpunkt att ytterligare begränsa möjligheterna till transport av vatten .
Detta skulle utgöra ett problem för de länder där vattenreserverna är ojämnt fördelade .
Ekologiskt hållbara transporter av vatten får inte begränsas genom unionens rättsakter .
Verksamheten skall givetvis också i fortsättningen vara reglerad och kräva tillstånd , men samma regler lämpar sig inte för till exempel Finland och Grekland som lider av torka .
Herr talman , fru kommissionär !
Vattnet är något naturligt och livsnödvändigt , och det är vår plikt att skydda det .
Jag anser det nödvändigt att det finns ett ramdirektiv för vattenpolitiken i Europeiska unionen , som kan bli det viktigaste rättsliga instrumentet för att förbättra vattenreservernas kvalitet och hantera dem på rätt sätt , och jag vill berömma föredraganden för hennes ansträngningar att ta itu med detta besvärliga problem och ta hänsyn till alla dess olika aspekter .
Jag måste emellertid påpeka att det i fråga om vatten finns skillnader mellan länderna i norr och länderna i söder , och därför kan man inte lösa vattenproblemen på samma sätt .
Det finns i Europa områden med strukturell vattenbrist , och detta måste man ta hänsyn till i direktivet .
Under de senaste åren har Medelhavsländerna , på grund av klimatförändringen , drabbats av allvarliga problem både i fråga om torka och i fråga om översvämningar .
Herr talman !
Jag stöder den gemensamma ståndpunkten , men jag accepterar också ganska många av de framlagda ändringsförslag som syftar till att förbättra den gemensamma ståndpunkten .
Däremot kan jag inte acceptera vissa andra ändringsförslag , t.ex. i fråga om prissättningen på vatten , med tanke på att en stor del av vattenanvändarna i vårt land är jordbrukare .
De ändringsförslag som vill förbjuda överföring av vatten mellan olika vattenreserver skulle leda till vattenbrist i många områden i mitt land .
Frågan om att få bort de skadliga ämnena måste vi hantera på ett mera realistiskt sätt , om vi skall lyckas .
Beträffande tiden för genomförande av direktivet måste man ta hänsyn till att det finns länder där infrastrukturen är sådan att det krävs både tid och avsevärda resurser för att genomföra direktivet .
Även efter dessa påpekanden , herr talman , anser jag att det gemensamma målet kvarstår , ett hållbart utnyttjande av vattenresurserna .
Herr talman , fru kommissionär !
Åtgärderna i föreliggande direktiv räcker allt ifrån iordningställande av planer för vattenförvaltning , omfattande information och rätt till utfrågning , intensivt samarbete mellan medlemsstaterna ända till bekämpning av vattenföroreningar som sker på grund av enskilda skadliga ämnen .
Och när man vet hur många år denna kammare har försökt att få ett sådant ramdirektiv , då gläder det mig att jag får vara med i dag , och jag vill gratulera Lienemann till att hon är den lyckliga som får lägga fram detta betänkande .
Men det är för mig mycket , mycket viktigt att också fastslå något som för många människor egentligen är självklart .
Trots detta vill jag betona följande : Detta direktiv erbjuder inte någon rättslig grund , hur den än ser ut , för att gentemot någon medlemsstats vilja leda bort vatten från dess område .
Och för att än en gång bekräfta detta har jag - tacknämligt nog med stort godkännande från PPE - lämnat in ett ändringsförslag , och det skulle glädja mig mycket om kammaren i morgon kunde rösta för mitt ändringsförslag .
Det handlar om ett klargörande att vattnet - och det har påpekats flera gånger i dag - inte är någon vanlig handelsvara , utan en tillgång som tillhör befolkningen i respektive medlemsstat i Europeiska unionen , och som måste skyddas och behandlas på lämpligt sätt .
Jag vet , och föregående talare har betonat det , att det finns stater i Europeiska unionen som har problem med vattnet .
Jag tror att vi i alla länder har möjlighet att behandla vattnet ännu bättre , och att se till att det används på ett ännu renligare sätt .
Inget land kan undantas från detta .
Men först när varje land har gjort en maximal ansträngning för att bevara sina vattenresurser , när allt verkligen har skett i det egna landet , först då , tror jag , bör det vara nödvändigt att tänka över ett solidariskt vattenutnyttjande .
Herr talman , fru kommissionär !
Det borde egentligen vara en anledning att glädjas att den andra behandlingen av detta direktiv redan är avslutad .
Ändå måste jag säga att jag inte känner någon glädje , för jag ser det som ett direktiv utan några större kvaliteter , som kommer att orsaka många problem och som har många brister .
Till att börja med kan jag säga att det är ett direktiv som är alldeles för tufft och förenklande , begränsande .
Tidigare direktiv på vattenområdet har sällan efterlevts och regeringarna och kommissionen har vid flera tillfällen undlåtit att kräva den disciplin som de borde , även om det är obehagligt .
Det är inte fråga om att man måste förfoga över mycket strängare regler , för problemen handlar många gånger om förvaltning , om att utöva sina befogenheter och inte till den lagstiftande makten överföra de omfattande problemen med vattensystemet , vars komplikationer vi alla är medvetna om .
Man har upprättat ett begränsande direktiv ; man kan inte låta det samma gälla för länder med segelbara floder som för länder där det råder brist på vatten , och där stora sprickor uppstår i marken på grund av vattenbrist och där det är 55º eller 60º i solen .
Jag säger detta , för bollen skall inte behöva ligga hos oss , utan bollen ligger hos regeringarna och kommissionen .
Likaså är den skadegörelse och de tragedier som äger rum , i Rumänien till exempel , inte problem som angår den lagstiftande utan den verkställande makten och regeringarna .
Det är dessutom inte ett solidariskt direktiv , för det bortser från de stora områdena , klimatskillnader , ökenområden , karga områden .
Det har upprättats med gemensamma kriterier som grund .
På området för överföring av vatten är det samma sak .
Att tala om överföring av vatten innebär att tala om fördelning av rikedom , av solidaritet mellan folk och mellan länder , för marken är tyvärr inte perfekt och vissa områden har mindre och andra har mer .
Slutligen ställer jag mig starkt kritisk till att direktivet inte åtföljs av en effektstudie .
Det är enkelt för oss att kräva av andra att de utvärderar effekterna men , vad miljön beträffar , bör vi kräva det av oss själva , med tanke på hur många människor , hur många jordbrukare som ruineras om de måste stå för kostnaderna .
Det har gjorts någon studie som inte ens har blivit läst , och jag anser att vi som god politisk tillämpning bör fastställa ett genomförande av miljöstudier ; i annat fall skapar vi doktrin .
Herr talman !
Genom sammanslagningen av nuvarande direktiv upprättas genom detta ramdirektiv den grundläggande principen för en hållbar vattenpolitik i Europeiska unionen .
Det är ett regelverk för att skydda och förvalta vårt vatten - ytvatten , grundvatten , övergångs- och kustvatten - genom att inrätta flodvattendistrikt på nationell och i vårt fall i Irland , på gränsövergångsnivå .
Irland stöder mycket den gemensamma ståndpunkten och många av Europaparlamentets ändringsförslag .
En period på 25 år för lagstiftning exempelvis är knappast godtagbart .
Vi har inga problem med principen " förorenaren skall betala " i förbindelse med omkostnadstäckning för vattennyttjande i fråga om industri- , handels- och jordbrukssektorn .
Jag har dock en bestämd åsikt att eftersom vatten är liv och tillgång till rent vatten en grundläggande mänsklig rättighet måste detta direktiv möjliggöra en gratis basförsörjning av hushållsvatten , en tilldelning per hushåll för dricksvatten , matlagning och sanitära ändamål .
Vi måste naturligtvis betala för slösaktig och överflödig användning i hushåll och omkostnadstäckningen kan balanseras i enlighet därmed .
Införandet av vattenmätare betraktas med stor misstänksamhet i Irland där vi inte har haft några avgifter för hushåll och följaktligen inga mätare sedan 1977 .
Mätare kan betraktas som ett mycket viktig verktyg för vattenförvaltningen av de nya flodvattendistrikten för att få bort vattenslöseri och för att kunna planera ordentligt för framtida behov .
Hela syftet med detta direktiv är att främja ett hållbart vattenutnyttjande i EU .
Vatten är en knapp och värdefull naturresurs .
I bästa fall skulle jag vilja att ändringsförslag 45 bortfaller i morgon så att den gemensamma ståndpunkten om artikel 9 skall gälla om vattenavgifter .
Det skulle ge möjlighet till subsidiaritet i fråga om kostnadspolicy för vattenavgifter där varje medlemsstat utformar sitt egen program så länge som detta direktiv om stimulansåtgärder för hållbart och effektivt vattenutnyttjande är fullständigt säkrade .
Om ändringsförslag 45 inte bortfaller skall jag var tvungen att lägga fram ett muntligt ändringsförslag i morgon för att säkerställa att medlemsstater får bevilja undantag till bestämmelserna i denna artikel och därmed göra det möjligt med en basvattenförbrukning för hushållsändamål innan avgifter debiteras för omkostnadstäckning .
All lagstiftning måste kunna verkställas och vara grundad på den allmänna principen om politiskt godkännande .
Jag anser att tillgång till rent dricksvatten utan avgifter är en grundläggande mänsklig rättighet i industriländerna liksom i utvecklingsländerna .
Herr talman , fru kommissionär , mina damer och herrar !
Nu när vi har kommit så här långt i debatten vill jag framhäva några aspekter som jag , från ett land i söder , ur agronomisk synvinkel anser vara av stor betydelse i detta direktiv .
Till exempel frågan om kostnaderna och frågan om överföring av vatten mellan magasin .
Vad beträffar kostnaderna , skulle jag vilja att vi specificerar vilka kostnader vi talar om .
Talar vi om resursernas fördelning och ursprung ?
Talar vi om distributionsnätens kvalitet ?
Talar vi om vilken typ av insatser som krävs för att de skall ge effekt ?
Eller talar vi om stora vattenbyggnadsarbeten och vattendammar ?
Summan av dessa kostnader som drabbar jordbrukssektorn skulle då bli gräsligt hög .
Vad beträffar överledningen av vatten kan det beskrivas som en överföring av ytvatten mellan de olika länderna .
Känner kommissionären till att vi vårt land har ett av de äldsta systemen för överledning av vatten i Europa ?
Sådana fanns för mycket länge sedan : redan på romarnas tid fanns de , men då var de mindre .
En av de viktigaste överledningarna - överledningen Tajo-Segura- , som har varit i drift i många år , i närmare 30 år , rymmer 658 hektometer3 / år .
Den största överförda mängden på ett år har varit 453 och genomsnittet under 20 år ligger på drygt tvåhundra .
Man kan inte anklaga oss för dålig förvaltning .
Känner kommissionären till att av dessa 263 hektometer3 är 25 avsatta till bevattning av västra Levante , 30 till försörjning av området Júcar , 7 till försörjning i den södra delen av Júcar och resten , i Segura , till lika stora delar försörjning och bevattning ?
Inte heller vi förvaltar detta på ett dåligt sätt .
Man kan inte förbjuda oss att göra överledningar när det är avgörande för vår ekonomi och för utvecklingen i våra områden .
Jag går inte in på frågan om kvalitet och de bästa tillgängliga metoderna , för jag tror att vi kommer att få förhandla om detta direktiv igen .
Men tänk på en sak : i det pluralistiska Europa som vi i solidaritet skapar måste vi eftersträva pluralistiska lösningar , inte unika lösningar .
Därför vädjar jag till förnuftet i kommissionen , i rådet och i denna församling , så att man vid omröstningen inte eftersträvar en enhetlighet mellan de olika europeiska länderna i frågor där subsidiariteten bör få råda .
Fru kommissionär : Andalusien är inte Lappland . .
Herr talman , ärade ledamöter !
Jag vill förstås börja med att tacka miljöutskottet och framför allt föredragande Lienemann för det ambitiösa och konstruktiva arbete som hon har lagt ned på detta ramdirektiv om vatten .
Vatten är en av våra viktigaste naturresurser , vilket många talare redan har sagt .
En ambitiös och välbalanserad europeisk politik på vattenområdet är en viktig del när det gäller att garantera en hållbar utveckling för Europa .
Vatten är också en av de frågor som jag kommer att ägna särskild uppmärksamhet åt under min mandattid .
Jag är glad för den anda av samförstånd som genomsyrar de ändringsförslag som har lagts fram för parlamentet .
Många av dem bygger på de mycket konstruktiva , informella diskussioner som fördes mellan parlamentet och rådet i samband med den första behandlingen .
De flesta av de ändringar som parlamentet föreslår bidrar till att förbättra texten och göra den mer ambitiös .
Kommissionen kan godta 72 av de 108 ändringsförslagen , antingen helt , delvis eller i princip .
Många av de ändringsförslag som parlamentet har lagt fram visar att en förlikning kommer att bli nödvändig .
Jag uppmanar därför parlamentet att med tanke på dessa kommande förhandlingar rösta för ett ambitiöst ställningstagande .
Först skulle jag vilja nämna några av mina viktigaste argument .
Vi har i dag möjlighet att sätta i verket de åtaganden som vi har gjort enligt Ospar-konventionen .
Hellre än att göra dessa målsättningar rättsligt bindande , måste vi se till deras politiska natur .
Detta reflekteras också i flera av parlamentets ändringsförslag .
Vad gäller vattenavgifter kommer detta direktiv att forma Europas vattenpolitik för de kommande tre årtiondena .
Det är vår skyldighet att redan i dag se till att detta direktiv ger de rätta incitamenten , de rätta drivkrafterna , för en effektiv avgiftsstruktur och prissättning som förbättrar vår miljö på ett kostnadseffektivt sätt .
Det låter bra att vatten skall vara en mänsklig rättighet och borde vara gratis .
Men vatten är inte gratis - lika litet som bostäder eller mat är gratis .
Det är först med effektiva styrinstrument som vi kan få en bättre hantering och en bättre hushållning med vatten .
Jag vill också tillägga att jag stöder en snävare tidsplan och förtydligande av mål och av undantagskriterier vad gäller grundvatten och vatten som är kraftigt modifierade av mänskliga aktiviteter samt att jag stöder det uttryckliga omnämnandet av radioaktiva ämnen .
Flera talare har under debatten påpekat hur viktigt det är med information och samråd med allmänheten .
Jag vill bara ytterligare understryka detta .
Det är helt avgörande att vi involverar allmänheten genom en bra information och genom ett samrådsförfarande .
Detta är också uttryckt i skäl 14 .
Låt mig också säga till Bowe att han såväl som min skotske medarbetare kan fortsätta att med gott samvete då och då smaka något glas skotsk whisky !
Vi har inte bedömt det vara nödvändigt att från kommissionens sida reglera det mycket begränsade uttaget av vatten för whiskyproduktion .
Låt mig nu få kommentera några av områdena litet mer i detalj .
Att begränsa utsläppen av farliga ämnen i våra vatten måste vara en av de viktigaste målsättningarna .
Jag är glad över att se att parlamentets ändringsförslag har koncentrerats på detta .
Kommissionen stöder helt förslaget att föra in Ospar-konventionens åtaganden i texten .
Vi måste dock hålla oss till deras exakta innebörd och räckvidd .
Som jag sade är målet och tidsplanen för Ospar främst ett politiskt åtagande .
Det skulle inte vara i överensstämmelse med detta att införa en rättsligt bindande tidsplan .
Det måste dock säkerställas att medlemsstaterna och gemenskapen tvingas vidta åtgärder för att uppnå dessa mål och följa tidsplanerna .
Jag välkomnar därför ändringsförslagen 6 , 10 , 14 , 24 , 58 , 60 och 88 .
Kommissionen kan däremot inte godta ändringsförslag 19 , där farliga ämnen definieras på ett annat sätt än i Ospar .
I kommissionens förslag införs ett tydligt förfarande för urval av ämnen , och därför behövs inte någon definition .
Även om jag också håller med om innebörden i ändringsförslag 79 och 106 , så går de utöver åtagandena i Ospar .
Jag kan därför inte godta dessa ändringsförslag .
Kommissionen kan också i princip godta ändringsförslag 60 , enligt vilket det krävs en tidsplan för kommissionens förslag om att begränsa utsläpp av prioriterade ämnen .
Ändringsförslag 59 inför krav på att förteckningen över prioriterade ämnen fortlöpande skall ses över .
Detta skulle medföra rättslig osäkerhet angående förteckningens status och kan därför inte godtas .
Begäran i ändringsförslag 60 och 93 om en målförteckning och en förteckning över ämnen , för vilka det inte finns tillräckliga data kan inte godtas .
Sådana förteckningar skulle få en oklar rättslig status och passar inte ihop med förfarandena för att anta förteckningen över prioriterade ämnen .
I detta sammanhang vill jag betona att Ospar-konventionen inte på något sätt förändrar den existerande gemenskapslagstiftningen vad gäller nitrat från jordbrukssektorn .
Nitratdirektivet kommer därför inte att påverkas av detta ramdirektiv .
Jag uppskattar att parlamentet visat sig vara flexibelt i den mycket känsliga och svåra frågan om att ta ut avgifter för vattentjänster .
Jag kan helhjärtat stödja kravet på att priset på vatten skall läggas på en nivå som innebär att det skapas incitament att använda vattenresurserna på ett hållbart sätt .
Jag stöder också kravet på ett lämpligt bidrag från varje sektor för att täcka de egna kostnaderna .
Jag kan därför delvis och i princip godta ändringsförslagen 43-46 samt ändringsförslag 85 .
Jag anser att vi behöver rättsligt bindande krav på att de finansiella kostnaderna för vattentjänster skall täckas av varje ekonomisk sektor .
Detta utgör ett tydligt mål i förhållande till vilket framsteg kan mätas .
Jag stöder därför den övergripande inriktningen i ändringsförslag 105 , som är i linje med kommissionens ursprungliga förslag .
Jag stöder också en successiv utveckling i riktning mot täckning av miljö- och resurskostnader .
Vi är medvetna om att priset på vatten och vattentjänster är en komplicerad fråga och att hänsyn måste tas inte bara till miljömål , utan även till sociala och ekonomiska mål .
Detta får dock inte vara en ursäkt för att subventionera förorenande och ineffektiva ekonomiska sektorer .
Vi har för avsikt att inom kort utfärda ett meddelande från kommissionen i just denna fråga .
Jag håller med parlamentet om att man avsevärt måste korta ned den tidsperiod för genomförandet på 16 år som anges i den gemensamma ståndpunkten .
Samma sak gäller även möjligheten som ges att förlänga genomförandet med ytterligare 18 år .
Ändringsförslag 28 som innebär att den tredje förlängningsperioden stryks är ett viktigt steg i rätt riktning .
Detta förslag kan därför godtas .
En period på tio år som föreslås bland annat i ändringsförslagen 24 och 26 är å andra sidan för kort .
Jag anser att man bör överväga att låta den övergripande definitionen av förslagets krav omfatta en uttrycklig och strikt bestämmelse om att undvika försämringar .
Förslaget måste också omfatta skärpta kriterier för förlängning av tidsfrister som gäller kraftigt modifierade eller konstgjorda vattenförekomster och för fastställande av lägre miljömål .
Detta gäller ändringsförslagen 6 , 24 , 25 , 27 , 30 , 31 , 32 , 33 , 34 , 78 , 80 , 102 och 104 .
Dessa ändringsförslag kan till väsentlig del godtas och kommer att stödjas för att en övergripande lösning skall kunna nås .
Kraven i ändringsförslag 27 och 29 , dvs , att kommissionen skall godkänna varje förlängning , skulle vara att gå för långt och kan inte godtas .
Ett annat viktigt område är skyddet av grundvattnet .
Vi behöver både en utgångspunkt och ett slutgiltigt mål för att vända den uppåtgående föroreningstrenden .
Vi behöver också strängare kriterier för tolkning av övervakningsresultaten .
De väsentligaste delarna av parlamentets ändringsförslag 25 och 73 kan därför godtas i princip .
Den nya definitionen i ändringsförslag 72 är dock för strikt och kan inte tillämpas i detta syfte .
Jag skulle föreslå att ändringsförslag 92 införlivas i en bredare lösning .
I ändringsförslag 71 tas inte hänsyn till årtidsvariationer och årliga förändringar i grundvattennivån .
Förslaget kan därför inte godtas .
Kommissionen anser det vara orealistiskt och onödigt att fastställa standarder genom vilka det säkerställs att den minst intensiva vattenreningen räcker till för att uppnå dricksvattenkvalitet av ytvatten .
I stället föredrar vi ett tillägg till de åtgärder som krävs enligt artikel 11 för att främja verksamhet på detta område .
Den goda status som krävs enligt detta förslag bör säkerställa att kravet på ytvatten av god kvalitet uppfylls .
Denna del av ändringsförslag 41 kan därför inte godtas .
Kommissionen uppskattar parlamentets insatser för att säkerställa att det så kallade kombinerade tillvägagångssättet ges en central roll .
Genom ändringsförslagen 22 och 47 definieras detta tillvägagångssätt och dess räckvidd , vilket kommissionen i princip kan godta .
För att uppnå största möjliga rättsliga tydlighet och proportionalitet vill vi dock formulera om ändringsförslag 47 och lägga till en de minimis-bestämmelse .
Överföring av vatten omfattas redan av kontroller , men ett uttryckligt omnämnande gör texten tydligare .
Denna del av ändringsförslag 49 och 87 kan således godtas .
Det är dock inte nödvändigt att fastställa som villkor att alla åtgärder för att styra efterfrågan vidtagits .
Förslaget fastställer redan att uttag av vatten måste ske i enlighet med de ekologiska behoven i ett avrinningsområde .
Denna del av ändringsförslag 49 och 87 kan därför inte godtas .
Kommissionen godtar ändringsförslag 76 som innebär att radioaktiva ämnen uttryckligen tas med i förslaget .
Sammanfattningsvis kan kommissionen godta 72 ändringsförslag helt , delvis eller i princip .
Följande ändringsförslag kan inte godtas : 1 , 4 , 9 , 11 , 13 , 15 , 19 , 23 , 39 , 40 , 51 , 59 , 61 , 64 , 66 , 70 , 71 , 71 , 72 , 74 , 77 , 79 , 81 , 83 , 87 , 89 , 90 , 91 , 95 , 97 , 98 , 100 , 101 , 103 , 106 , 107 .
Avslutningsvis vill jag säga att jag välkomnar de ansträngningar som parlamentet har gjort för att försöka lösa de frågor som rådet har en annan uppfattning om .
Viktiga framsteg har gjorts och den konstruktiva tonen i diskussionerna skapar ett bra arbetsklimat för framtida förhandlingar .
Ett antal hinder återstår , men jag är övertygad om att vi i takt med att lagstiftningsarbetet går vidare kommer att uppnå vårt gemensamma mål om att skapa en vattenpolitik , som vi kan vara stolta över .
Ett bestämt ställningstagande från parlamentet sida kommer att vara ett viktigt bidrag till en ambitiös , europeisk vattenpolitik för de närmaste tre decennierna .
( Applåder ) Jag skulle vilja höra kommissionärens åsikt om ändringsförslag 45 .
Jag kanske missade den i den förteckning som delades ut . .
( EN ) Jag godtar det .
Tack för det , fru Wallström .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.30 .
 
Finansiellt instrument för miljön ( Life ) Nästa punkt på föredragningslistan är andrabehandlingsrekommendation ( A5-0014 / 2000 ) från utskottet för miljö , folkhälsa och konsumentfrågor om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om det finansiella instrumentet för miljön ( Life ) ( Föredragande : Marie-Noëlle Lienemann ) . .
( FR ) Herr talman , vi fick redan tillfälle vid första behandlingen att granska betänkandet och jag trodde mig förstå i utskottet att det fanns ett stort samförstånd i församlingen .
Life är den enda budgetposten i gemenskapens budget för en direkt insats på miljöområdet och vi måste konstatera att den inte är i nivå med våra ambitioner eftersom de summor som den får har stagnerat i åratal : trots utvidgningen som redan hade ägt rum då vi förnyade det första Life-programmet för att gå över till det andra , trots utvidgningen hade anslagen bibehållits .
Och sedan ser vi att regioner , olika aktörer , företag , sammanslutningar mer och mer lämnar in Life-projekt , såväl till Life " natur " som Life " miljö " , och att dessa projekt har mycket god kvalitet och efter en teknisk granskning av samtliga behöriga kommittéer är alla överens om att säga att de skulle förtjäna stöd av Europeiska unionen och vi lyckas ändå inte finansiera dem i brist på budgetanslag .
Man måste också påminna om att denna budget är föremål för en exceptionell anslagsförbrukning i gemenskapens budget .
Vi har således här uppenbarligen ett redskap som är väl anpassat för den politik som vi vill genomföra .
Och jag vill särskilt framhålla avdelning Life " natur " .
Vi vet att i Europeiska unionen möter en hel rad direktiv rörande " Habitat " direktivet och direktivet om " Flyttfåglar " tillämpningssvårigheter : vi borde kunna ledsaga Life " natur " med de politiska åtgärder som visar på genomförbarhet , berättigande samt kapacitet att genomföra målsättningarna i direktiven .
Och i brist på anslag förlorar vi denna legitimitet låter tanken utvecklas att våra europeiska direktiv inte är rimliga och tillämpliga .
De debatter som sålunda äger rum i dag koncentreras på två stora ämnen : i första hand , kommittéförfarandet , den eviga debatten i kammaren , men parlamentet ville vidta politiska åtgärder som snarare slutar med förvaltningskommittéer och samrådskommittéer som ger en viss flexibilitet åt kommissionen och ger inte alltför mycket kapacitet åt rådet att låsa och göra gällande , skulle jag säga , regeringsfilosofin jämfört med gemenskapsfilosofin som vi står som garant för här i Europaparlamentet .
Men debatterna om kommittéförfarandet har vi med anledning av de flesta av Europeiska unionens finansprogram och finansredskap .
Jag skulle säga , verkar det som , - och de kontakter som vi har kunnat få tenderar att visa det - att , säger jag , närmanden av synpunkter om kommittéförfarandet förvisso är lättare än budgetnärmanden .
Jag vill påminna om att parlamentet kräver anslag på 850 miljoner ecu , vilket inte är enormt i gemenskapsbudgeten , och att de aktuella förslagen ligger på 613 miljoner ecu .
Det tycks mig i varje fall som att åtminstone mot slutet av tillämpningen av Life skulle det finnas möjlighet för unionen att göra en betydande budgetgest till förmån för miljön .
Låt mig sluta med frågan om våra institutioners sätt att fungera .
De uttalanden jag hör nu är : " Vi måste absolut lyckas avsluta snabbt nu . "
I klartext , i parlamentet drar ni ner era anspråk , i synnerhet era budgetanspråk !
För om vi inte lyckas snabbt inom ramen för medbeslutande att fastställa ramen för Life-förordningen skall vi försenas i genomförandet för år 2000 och visserligen väntar de icke-statliga organisationerna , aktörerna i terrängen , på våra anslag .
Jag skulle emellertid vilja påminna om att rådet förfogar över en mycket lång tid för att göra sig en idé och att det inger sina förslag några månader före den ödesbestämda tidsfristens utgång .
Vi för vår del , vi är bundna av texterna : maximalt fyra månader .
Vi håller våra tidsfrister och efteråt säger man : " Vänta !
Om ni vill vara förnuftiga , får ni acceptera vår ståndpunkt , eftersom det inte finns någon tid i medbeslutandeförfarandet " .
Jag tror att vårt parlament ofta protesterar mot denna metod som inte ifrågasätter någon särskild person i rådet och jag skulle absolut inte vilja att det portugisiska ordförandeskapet känner sig skyldig till detta tillstånd eftersom det i verkligheten är litet av en tradition som rådet uppehåller i tiden .
Men jag skulle vilja insistera på att budgetfrågan är central för denna miljöfråga och att parlamentet inte kan ge efter för den utpressning som skulle tvinga det att vara den enda förnuftiga i denna fråga .
Jag hoppas således att våra kolleger kommer att stödja oss i förlikningen - men omröstningarna har alltid varit mycket överensstämmande i den dimensionen - men också att rådet och kommissionen kommer att lyssna på oss och att vi kommer var och en att ta ett steg mot varandra .
Herr talman , ärade kollegor !
Det är sant att vi är öppet oense vad gäller en del av de alternativ som rådet och kommissionen har valt .
Detta har jag dock en möjlighet att ta upp litet längre fram .
Samma sanning manar mig emellertid att börja med att säga att den här regleringen är bättre än den som hänför sig till Life I och Life II .
Först och främst för att Life blev striktare , öppnare och mera rationell tack vare det grundläggande förslaget .
För det andra för att man i den gemensamma ståndpunkten integrerar några fundamentala synpunkter , definierade av Europaparlamentet vid den första behandlingen , nämligen att sysselsättningsskapande åtgärder skall vara en faktor att ha i åtanke när kandidatprojekten väljs samt att en produkts globala påverkan från tillverkning till återvinning och eliminering skall minskas och vara ett av de mål man vill nå med Life miljö .
För det tredje är vi mycket positivt inställda till det faktum att man i den gemensamma ståndpunkten för första gången tog med värdestegring och territoriella bestämmelser för kustområden som en av de frågor som Life miljö skall prioritera .
Herr talman , ärade kollegor , trots alla dessa dygder så fallerar man när man inte låter Life III reglera det som är så uppenbart och viktigt för effekten av ett finansiellt instrument : dess budget .
Genom att stå fast vid sitt förslag om 613 miljoner euror som referensbelopp för perioden 2000-2004 och genom att förhindra Europaparlamentets förslag om 850 miljoner euror står kommissionen och rådet i begrepp att fatta ett beslut som enligt vår mening inte grundar sig på samma omdömesförmåga och samma rättvisekriterier som man så omsorgsfullt har introducerat i andra förordnanden i Life III .
Kommissionen och rådet skall veta att vi från vår sida inte kommer att ge oss förrän Life har försetts med den budget den förtjänar och som på bästa sätt kan borga för att de miljöresultat man vill uppnå med ett sådant instrument verkligen uppnås .
Vi rättfärdigar vårt val med fyra mycket enkla argument .
För det första så är Life det enda direkta finansiella instrument som finns för att gynna miljöpolitiken inom Europeiska unionen .
Det finns inget annat .
För det andra så är Life ett instrument som man har åstadkommit goda resultat med , som man har utvecklat metoder och ny teknik med som till stora delar har förverkligats .
För det tredje så har budgeten för Life reellt sett minskat och den har inte följt den enorma dynamik och kreativitet som man velat .
För det fjärde så har parlamentet , tack vare den betydelse som tillskrivs Life , i sin årliga budget höjt sina anslag till det här programmet , vilket gör att ett godkännande av det förslag som rådet och kommissionen tar i försvar skulle innebära en oacceptabel vändning av den tendensen .
Vi är dock inte bara oroade över budgetfrågan .
De klimatologiska förändringarna och vattenpolitiken är frågor som de europeiska medborgarna oroar sig mycket för och som förtjänar kammarens odelade uppmärksamhet .
Därför är det viktigt för oss att våra ändringsförslag 5 och 6 godkänns , där man försöker definiera en hållbar förvaltning av käll- och ytvatten samt en reducering av växthusgaser som mål att nå med Life miljö .
Ett sista ord för att tacka ledamot Lienemann för hennes betänkande , samtidigt som jag passar på att berätta att vi kommer att rösta för ändringsförslagen om kommittéförfarandet även om vi hade föredragit , som det så påtagligt kom fram i utskottet för miljö , att Life hade åtföljts av en rådgivande kommitté , så vill vi inte bidra till att rådets förslag går igenom , ett förslag som uppriktigt sagt är betydligt sämre .
Herr talman !
Fru kommissionär !
Fru kommissionär , ni utövar med all rätt press på de medlemsstater som inte har genomfört direktivet om livsmiljöer samt vilda djur och växter , också på den medlemsstat som jag kommer från .
Detta med all rätt , eftersom kraven på våra naturliga livsrum finns kvar och vi äntligen måste genomföra dessa Natura-2000-områden .
Men när detta sker , då har vi naturligtvis ett enormt behov av Life-Natura-pengar , eftersom vi i dessa områden , som då äntligen legitimeras , naturligtvis också måste finansiera åtgärder för att bibehålla dem , och detta i en situation där vi inte en gång kan stabilisera det som vi har uppnått med Life I och II .
Med tanke på denna situation , att områden för att bevara livsmiljöer samt vilda djur och växter nu måste tvingas fram , behöver vi entydigt också mer pengar för Life .
Här vänder jag mig också till rådet : Rådet är världsmästare när det gäller att besluta om utgifter just när det gäller utrikespolitiken , som vi sedan på något sätt måste finansiera med vår budget .
Jag kan bara nämna hjälpen till Bosnien - där gör vi nedskärningar på alla möjliga områden .
Här däremot vägrar rådet att i ett längre perspektiv utöka Life-budgeten med belopp som ändå är skrattretande i förhållande till den totala budgeten , på ett område där det dock handlar om vår hållbara utveckling .
Det kan jag inte på något sätt förstå , och jag ber alla kolleger eftertryckligen att stödja kollegan Lienemanns förslag om en höjning till 850 miljoner euro .
Herr talman , kära kolleger !
Life är i själva verket Europeiska unionens viktigaste instrumentet , det enda finansiella instrumentet , som enbart är ägnat åt miljö .
Därmed är det sagt att detta redskap bör vara i nivå med våra ambitioner , ambitioner som har ett pris , naturligtvis .
Den grundläggande diskussionspunkten med rådet kommer självklart att vara det anslag som Life III bör ha .
I den gemensamma ståndpunkten planerades ett finansiellt totalanslag på 613 miljoner euro för perioden 2000-2004 , det räcker inte .
Den liberala gruppen är positiv till en ökning av beloppet till 850 miljoner euro .
Vi stöder således Lienemanns ändringsförslag som noterar att anslaget för Life inte ökades vid den senaste utvidgningen av unionen , för att ändå inte tala om nästa tåg med nyanlända .
De summor som vi begär är inte ett Himalaya med onödiga utgifter .
Tvärtom de förblir anspråkslösa i förhållande till de behov som skall täckas .
En droppe i havet - skulle jag säga - jämfört med Europas strukturpolitik .
Miljön förblir den fattiga kusinen i den europeiska budgeten samtidigt som den framför allt utgör en investering .
En investering i naturresurser naturligtvis men också i sysselsättning , eftersom det har bevisats att en aktiv miljöpolitik skapade nya arbetstillfällen , beviset är i synnerhet den mycket stora framgången med Life : en framgång hos icke-statliga organisationer , företag , lokala myndigheter samt tredje land .
Nära en tredjedel av 8 500 mottagna efterfrågningar uppfyllde kraven och omkring 1 300 projekt samfinansierades mellan 1992 och 1998 .
En framgång som parlamentet vill se och ämnar se till att den fortsätter , vilket är skälet till att vi också stöder ändringsförslag 14 som drar upp den fjärde etappen under Life-projektets livstid .
När det är fråga om miljö , minskar investeringar och ambitioner och skall minska på lång sikt .
Det är priset för de kommande generationernas framtid .
Herr talman , fru kommissionär !
Jag kommer utan tvivel att upprepa vad mina kolleger sagt , men jag tror att vad beträffar rådet handlar det om att upprepa gång på gång vad vi tycker om Life .
Jag kommer således också att säga - såsom föredraganden redan har gjort så bra - att Life är det enda specifika finansiella instrumentet för införandet och genomförandet av Europeiska unionens politik på miljöområdet .
Detta instrument är absolut väsentligt eftersom det ger impulser till verkligt nydanande åtgärder till förmån för natur och miljö i Europa , vilket tas upp och förstärks av medlemsstaterna .
Detta finansiella instrument är för övrigt med vilja demokratiskt genom att det är lika tillgängligt för statliga organisationer som för icke-statliga organisationer .
Kära kolleger , därför ber jag er att inte rösta för de ändringsförslag som inte har förstått någonting om Lifes anda .
Life är direkt användbart av den europeiska medborgaren via sammanslutningar och för åtgärder av allmänt intresse .
Flera miljoner - jag sade miljoner - medlemmar i icke-statliga organisationer känner i Life unionens vilja att bygga upp en ambitiös politik till förmån för naturarvet .
Life är för övrigt ett grundläggande instrument för nätet Natura 2000 i Europa på vilket medlemsstaterna satsat , i enlighet med gemenskapsdirektiven om bevarande av livsmiljöer samt vilda djur och växter och om flyttfåglar , vilket gör det möjligt att införa skydd av platser av högt biologiskt värde i våra stater .
Jag skulle vilja säga att de som avböjer denna politik i sina stater bär ansvaret att bromsa naturskyddspolitiken i Europa .
Det är synd , eftersom alla vet i denna kammare att Life är ett otillräckligt finansiellt instrument för att genomföra de projekt som läggs fram av medlemsstaterna , varav många avslås i brist på finansiella medel .
Vi får inte glömma att Life bara får 100 miljoner euro per år , det vill säga knappt en promille av unionens budget .
Till påminnelse kan sägas att jordbruket , vars påverkan på miljön är reell får en budget på - vi vet alla - 37 miljarder euro .
I det sammanhanget anser min grupp att det är absolut nödvändigt att öka anslaget för Life och stöder reservationslöst Lienemanns förslag att öka budgeten till 850 miljoner euro , eftersom vi vet - jag tror att man måste säga det - hur stark förväntan är bland medborgarna i fråga om miljön och hur mager och oacceptabel kompromissen från rådet är rörande budgeten för Life , framför allt som Life-programmen har exceptionell verkställighet och har visat i vilken grad de gör det möjligt att framkalla nya miljömetoder .
De första projekten för hållbar utveckling är utan tvivel dessa projekt .
Herr talman , Europeiska unionens miljöprogram , som tilldelats avsevärda medel ( 613 miljoner euro ) ställer många frågor om ett gott utnyttjande av offentliga medel .
Ett finansiellt instrument av denna betydelse måste vara öppet och effektivt , vilket inte är fallet av följande skäl : dåligt definierade urvalskriterier , tvivelaktiga och åtgärder som kommit till utan samråd , icke offentliggjorda sammanfattningar , frånvaro av utvärderingspolitik .
Vi föreslår er således att ändra förordningen på följande sätt .
För det första , skall förvärv som görs med Life-medel endast förbehållas offentliga strukturer , även om förvaltningen av platserna anförtros efter anbudsinfordran åt sammanslutningar som auktoriserats för naturskydd .
Inköpens varaktighet är beroende av det , eftersom privaträttsliga sammanslutningar kan försvinna eller sälja vidare .
Det är filosofiskt chockerande och rättsligt bestridligt att 100 procent av offentliga pengar skall användas för att bygga upp privata fastighetstillgångar , till och med under miljöskyddets täckmantel .
För det andra , skall kriterier för stödberättigande och tilldelning av Life-medel fastställas för att undvika misstankar om kundgynnande och ostracism .
För det tredje , skall det i förväg krävas ett samråd med de berörda användarna och myndigheterna .
Till exempel , Life-natur i Frankrike , Grand-Lieu , som utarbetades utan något samråd ledde till en verklig ekologisk katastrof , eftersom slamborttagandet , som gjordes utan hänsyn till den franska vattenlagen , ledde till en betydande uppslamning av Acheneau , ett vattendrag uppströms , med förstörda fisklekplatser och utfyllda våtområden och så vidare .
Man flyttade nämligen slammet tre kilometer till en kostnad på sex miljoner franc , en bot som var värre än det onda , en förutsedd konsekvens som förebådades av alla aktörer på platsen .
Resultatet blev ett tvistemål och en kostnad för återställande som var högre än programbeloppet .
Det är vad vi vill undvika .
För det fjärde , skall det i uppföljningskommittén ingå företrädare för parlamentet och minst en ledamot per politisk grupp .
Att ledamöterna följer användningen av de röstade anslagen är väl legitimt ?
För det femte , skall årligen en vetenskaplig , teknisk och finansiell sammanfattning offentliggöras om de genomförda Life-åtgärderna .
För det sjätte , skall en seriös och regelbunden utvärdering av programmen ske .
För det sjunde skall dessa fonder kunna användas i händelse av miljökatastrof : till exempel , för trädplantering efter storm , återställande av naturområden efter oljeutsläpp , osv .
Fru föredragande , herr talman , här har ni nu detta förslag som är konkret , förnuftigt , lätt att genomföra , av den karaktären att det begränsar lokala konflikter och rättfärdigar en god användning av offentliga pengar och som vi föreslår före alla ökningar - plus 40 procent i alla fall ! - av budgetposten för Life .
( Applåder ) Herr talman , fru kommissionär , mina damer och herrar !
Jag vill börja med att gratulera Lienemann till det betänkande hon har upprättat och även kommissionen - varför inte - eftersom detta betänkande , detta ställningstagande , rent allmänt förbättrar de texter som är gällande .
Dessutom är systemet bättre och betänkandet är tydligare och mer genomblickbart .
Jag vill även gratulera kommissionstjänsten , till att utvärderingen , kontrollen och uppföljningen av programmet Life på ett förnuftigt sätt garanterar urvalet och genomförandet av projekten .
Däremot finns det några punkter jag vill ta upp .
För det första kontinuiteten som jag i princip inte ifrågasätter .
För det andra de finansiella anslagen .
Tyvärr är det endast 7,2 procent av de föreslagna projekten som finansieras .
Av de begärda 1 919 miljoner euro beviljas endast 784 miljoner euro i anslag .
I budgetplanen förekommer endast 613 miljoner euro till övriga länder och befogenheter .
Parlamentet har redan föreslagit 850 miljoner euro , men i dokumentet upprepas det första förslaget , 613 .
Fru kommissionär , miljötvånget växer på alla områden samtidigt som det enda finansiella instrumentet som endast är avsett för miljön minskar .
Är inte det en motsägelse ?
Begär vi av andra det vi inte är beredda att ge ?
Varför talar vi alla så mycket om miljön , när vi inte är beredda att tillsammans finansiera denna , utan i stället vill att den skall finansieras och bevaras av dem som bor där året om ?
Fru kommissionär , låt oss vara konsekventa .
Kostnaderna för att bevara den miljö som vi alla njuter av bör vara allas ansvar , och programmet Life är det enda finansiella instrumentet som endast är avsett för miljön med projekt som i regel brukar ha god verkan .
Herr talman !
Life är sedan 1992 gemenskapens främsta instrument för att stödja och utveckla miljöpolitiken såväl inom gemenskapen som i förbindelserna med tredje länder .
Med stöd av de senaste åtta årens erfarenheter försöker man att effektivisera miljöinsatserna i detta finansiella instruments tredje fas .
Viktiga inslag i den förordning vi skall rösta om är finansiering av insatser för att tillämpa , anpassa och utveckla gemenskapens politik på miljöområdet men också hänsynstagandet till miljöaspekter inom andra politikområden och strävan efter en hållbar utveckling .
I avsnittet Life-natur , som framför allt tar sikte på förverkligandet av naturnätverket 2000 , är det betydelsefullt att man anlägger ett mångnationellt perspektiv vid utarbetandet av internationella projekt och insatser , så att man undviker en uppsplittring av biotoperna , samtidigt som man ökar skyddet av den biologiska mångfalden .
I det andra avsnittet , Life-miljö , som framför allt gäller demonstrationsprojekt för de små och medelstora industriföretagen och organen för lokal självstyrelse , sägs det uttryckligen att miljöpolitiken måste införlivas i de övriga politikområdena .
När det gäller finansieringen av Life under de följande fem åren , instämmer jag i föredraganden Leinemanns förslag om en ökning från 613 miljoner euro till 850 .
Det ökade miljömedvetandet och hänsynstagandet till miljöaspekterna under de senaste åren får ingen effekt , om man inte kan få fram nödvändiga resurser för miljöskydd .
Vi kan heller inte vara likgiltiga för de växande problemen i unionens omvärld eller de akuta miljöproblemen i ansökarländerna .
Ett tydligt exempel är den giftkatastrof som nyligen inträffade i Donau och i en av dess bifloder .
Jag anser alltså att insatserna för ökat miljöskydd genom finansieringsinstrumentet Life är en garanti för att gemenskapens miljöpolitik skall lyckas och att de på ett betydelsefullt sätt hjälper gemenskapen i dess uppgift att skydda och förbättra miljön .
Herr talman !
Först av allt vill jag gratulera Lienemann till den starka känsla för miljöfrågorna som märks i de två betänkanden vi diskuterar i kväll .
Två minuter är verkligen inte tillräckligt för att avhandla ett så viktigt ämne .
Jag skall därför bara rikta en vädjan till kommissionären att hon tar med sig detta så ansenliga bagage .
Sedan fem år är jag ansvarig för miljöutskottet i en annan institution som , eftersom den har regional karaktär , verkligen inte har så vida vyer som detta parlament .
Miljösituationen är mycket , mycket allvarlig .
Liksom de kolleger som talat före mig skulle jag än en gång vilja uppehålla mig vid frågan om ekonomin och finansiering av projekt som , enligt min mening , alla borde ha offentlig karaktär .
Finansieringen : Fru kommissionär , 613 miljoner euro räcker inte .
Inte heller 850 miljoner euro räcker .
I slutet av augusti deltog jag vid ett möte med utskottet för miljö där man talade om 2 miljoner euro rent av , eller 4 000 miljarder lire , för att eliminera eller åtminstone minska nikotinproblemen .
Och ändå är miljön ett mycket allvarligare problem , mycket viktigare än rökningen .
Jag försäkrar er , fru kommissionär , att 850 miljoner euro - under förutsättning att dessa medel verkligen har avsatts - inte räcker för att i praktisk verklighet driva någon form av projekt .
På många håll har man anlagt parker , som enligt Life-programmet är av grundläggande betydelse .
Men parker som anläggs med knappa ekonomiska medel , utan skyltning , är ineffektiva och onödiga .
Därför uppmanar jag parlamentet och kommissionen att noga följa denna fråga . .
Herr talman , ärade ledamöter !
Ända sedan början av 1999 har det förts diskussioner mellan institutionerna om den föreslagna förordningen för en tredje etapp för instrumentet för miljön - Life .
Jag vill återigen tacka miljöutskottet och Lienemann för det goda och konstruktiva samarbete som vi har haft i detta ärende .
Som ett resultat av det kan jag bekräfta att kommissionen helt eller i princip godtar nio av de fjorton ändringsförslag som har antagits i miljöutskottet .
Kommissionen välkomnar framför allt ändringsförslagen 1 , 2 , 7 , 8 , 9 , 10 , 11 och 13 , som gäller kommittéförfarandena .
Parlamentet har i dessa fall helt beaktat de invändningar som kommissionen hade mot den gemensamma ståndpunkten .
Kommissionen kan i princip också godta ändringsförslag 4 , som dock bör föras in på ett annat ställe i texten .
När det gäller ändringsförslagen 5 och 6 vill jag betona att projekt för ett hållbart nyttjande av grundvatten och ytvatten samt projekt för minskning av luftföroreningar som bidrar till växthuseffekten i stor utsträckning omfattas av Life .
Kommissionen anser dock att man , om man anger detta separat , går emot det ursprungliga beslutet att koncentrera förslaget till några få prioriterade områden .
Det finns också en risk för överlappning med andra gemenskapsprogram som femte ramprogrammet för forskning , teknisk utveckling och demonstration .
Detta programs nyckelåtgärder - vattenkvalitet , morgondagens stad och innovativa produkter och processer - omfattar till viss del samma frågor .
När det gäller budgetfrågan är jag glad över det förtroende som miljöutskottet visat .
I ändringsförslag 12 begärs en större budget än den som anges i den gemensamma ståndpunkten .
Jag är också övertygad om att Life har stor potential .
Detta instrument skulle kunna finansiera bra projekt med ett högre belopp än det som anges i den föreslagna budgeten .
Det belopp som anges i ändringsförslag 12 är dock inte i enlighet med den budgetplan som fastställts på grundval av Agenda 2000 .
Låt mig också få foga in att om man höjer budgeten är det självklart att det också krävs mer av miljödirektoratet för att hantera ett ökat antal projekt .
Hänsyn måste också tas till andra program om vilka beslut skall fattas inom ramen för medbeslutandeförfarandet .
Kommissionen håller i detta skede fast vid det belopp som fastställts i den gemensamma ståndpunkten .
När det gäller ändringsförslag 3 , som vi inte godtog vid den första behandlingen , vill jag betona att varje program har sina egna mål , stödberättigande kostnader och ansökningsbestämmelser .
Det är därför meningslöst och ofta omöjligt att direkt överföra projekt från Life till andra instrument .
Om man för varje projekt skulle undersöka andra finansieringskällor , skulle det dessutom krävas mer resurser än vad som i dagsläget finns att tillgå .
Nu när kommissionen noga måste överväga vilka resurser som krävs för varje verksamhet är detta ett exempel på en icke central , men resurskrävande verksamhet som vi bör undvika .
Kommissionen kan inte heller godta ändringsförslag 14 , som står i strid med kommissionens initiativrätt .
Beträffande diskussionen om slutdatum vill jag säga att det slutdatum för att börja genomförandet av Life , den 31 mars år 2000 , som sattes i den gemensamma ståndpunkten nu måste flyttas fram .
Datum kommer att fastställas så fort denna förordning är antagen .
Avslutningsvis vill jag upprepa att jag är övertygad om att Life kommer att bli ett verkningsfullt instrument till stöd för utvecklingen och genomförandet av gemenskapens miljöpolitik .
Parlamentet har i stor utsträckning bidragit till att förbättra detta instrument .
Jag är övertygad om att ni delar min önskan om att förordningen skall kunna antas så snart som möjligt , speciellt med tanke på att det finns stora förväntningar i medlemsstaterna och i andra länder , inte minst bland kandidatländerna som nu ges möjlighet att delta i Life .
Tack för det , fru Wallström .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.30 .
 
Modernisering av social trygghet Nästa punkt på föredragningslistan är betänkande ( A5-0033 / 2000 ) av Andersson för utskottet för sysselsättning och socialfrågor om meddelandet från kommissionen -En samordnad strategi för att modernisera social trygghet ( KOM ( 1999 ) 347 - C5-0253 / 1999 - 1999 / 2182 ( COS ) ) . .
Herr talman !
Frågan om de sociala trygghetssystemen är en viktig fråga .
Detta är en naturlig följd av samarbetet inom EU .
Grunden är det monetära samarbetet , som sedan har följts upp av ett makroekonomiskt samarbete och ett samarbete om sysselsättningspolitiken .
Nu är det en naturlig följd att gå vidare med de sociala trygghetssystemen .
Dessa områden är ömsesidigt beroende av varandra .
Ekonomisk stabilitet är en grund för tillväxt och kan ge en hög sysselsättning .
Det ger också möjlighet att utveckla välfärden .
Det omvända förhållandet gäller emellertid också : en väl utvecklad politik när det gäller den sociala tryggheten kan bidra till hög sysselsättning och till en ökad tillväxt .
Social trygghet är med andra ord en produktiv faktor .
Det finns skillnader inom EU när det gäller de sociala trygghetssystemen .
Mycket av detta är historiskt betingat .
Nu har vi dock ett antal gemensamma utmaningar framför oss .
Det gäller exempelvis den demografiska utvecklingen som inte bara handlar om att antalet åldringar ökar , utan även om ett minskat barnafödande .
Arbetsmarknaden förändras också .
Kvinnor söker sig i allt större utsträckning ut på arbetsmarknaden .
En annan utmaning är den tekniska utvecklingen .
Dessa utmaningar måste vi möta gemensamt .
Kommissionens meddelande förordar ett ökat erfarenhetsutbyte samt att en högnivågrupp bildas och att benchmarking skall ske .
Dessutom skall rapporten om social trygghet ges ut årligen och granskas tillsammans med sysselsättningsrapporten .
Detta är bra , men det räcker inte .
Vi föreslår ett förfarande likt Luxemburgprocessen .
Det behövs tydliga riktlinjer och indikatorer , samtidigt som medlemsstaterna skall utforma metoderna i nationella handlingsplaner .
Vi skapar en gemensam modell , men bevarar subsidiariteten .
Denna sociala konvergens är en process som kommer att fortgå under lång tid .
Därför måste parlamentet involveras i arbetet - inte genom att ingå i högnivågruppen , men genom att företrädare för parlamentet kan följa arbetet i högnivågruppen och komma med förslag om hur processen skall bedrivas .
Kommissionens förslag är likt sysselsättningssamarbetet uppbyggt på fyra pelare .
Dessa är : att göra systemen sysselsättningsvänliga , att göra pensionssystemen långsiktigt hållbara , att främja social integration och att garantera en hållbar hälso- och sjukvård av hög kvalitet .
Allt detta är viktigt .
I vårt betänkande har vi särskilt pekat ut vikten av att bekämpa fattigdomen inom EU och att snarast möjligt finna indikatorer så att vi kommer framåt på detta område .
Jämställdheten har ingen egen pelare .
Det är mainstreaming som gäller .
Jämställdhetsaspekter skall därför återfinnas inom alla fyra pelarna .
Detta har vi tagit fasta på .
Vi lägger fram en mängd förslag , t.ex. om en övergång till individualiserade sociala trygghetssystem , att föräldraledighet skall kvalificera till förmåner i de sociala systemen , förbättrade möjligheter att förena familje- och arbetsliv , samt att den grundläggande ålderspensionen skall garantera en anständig levnadsnivå .
Dessa förslag gynnar framför allt kvinnor .
Parallellt med denna europeiska sociala konvergensstrategi krävs en konkret plan för lagstiftningsarbete på det sociala området samt förslag till ramavtal inom ramen för den sociala dialogen med en konkret tidsplan .
Vi förväntar oss att kommissionen presenterar detta i sitt förslag till socialt handlingsprogram .
Den sociala konvergensen är också nödvändig inför utvidgningen , dels för att stärka den sociala modellen , dels för att bekämpa riskerna med social dumpning .
Kommissionen bör överväga att ta fram ett särskilt handlingsprogram beträffande socialpolitiken i samband med utvidgningen .
Vi har i utskottet fört en konstruktiv diskussion .
Vi hade många ändringsförslag , men lyckades enas om ett betänkande .
Nu har de ändringsförslag som går till omröstning i plenum minskat till endast femton .
Detta tyder på att vi har en stor samsyn .
En del av dessa ändringsförslag återkommer från utskottsbehandlingen .
Dem kommer jag att avvisa .
Jag kommer också att avvisa de ändringsförlag som lagts fram av TDI-gruppen , eftersom jag inte tycker att dessa tillför betänkandet något .
Däremot kommer min grupp att bifalla ändringsförslag 14 från den liberala gruppen .
Detta förslag tycker jag är bra .
Visserligen liknar det ändringsförslag 1 , men ändringsförslag 14 är bättre .
Avslutningsvis vill jag säga : EU handlar inte bara om handelssamarbete .
EU handlar också om en union för sysselsättning och social rättvisa .
I skapandet av ett medborgarnas Europa spelar socialpolitiken en viktig roll .
Parlamentet vill med detta betänkande lämna sitt bidrag till en förstärkt social dimension i det europeiska samhället .
Vi hoppas att rådet och kommissionen tar detta bidrag på allvar och tar med det i den framtida socialpolitiken .
Toppmötet i Lissabon är ett utmärkt tillfälle att presentera en sådan strategi .
Herr talman , fru kommissionär , mina damer och herrar !
Ett långsiktigt bärkraftigt socialt trygghetssystem , där män och kvinnor på lika villkor har en trygghet som motsvarar deras särskilda livssituationer , är absolut nödvändigt för den sociala sammanhållningen och för stabiliteten i vårt samhälle .
Det ömsesidiga beroendet när det gäller ekonomin i sin helhet , sysselsättningspolitiken och den sociala tryggheten på den inre marknaden kräver här också gemensamma överläggningar på gemenskapsnivå .
Någon jämställdhet för män och kvinnor har inte uppnåtts varken inom arbetslivet eller i fråga om den sociala tryggheten .
Arbetslösheten är betydligt högre för kvinnor än för män .
Kvinnor har fortfarande sämre tillgång till yrken , och deras andel av besvärliga arbeten och deltidsarbeten är mycket högre .
Kvinnornas lönenivå ligger fortfarande långt under männens .
Det resulterar i en dålig social trygghet , eller fullständig brist på den , eftersom det enligt gällande system är det betalda arbetet som tjänar som grundval .
Många kvinnor åtnjuter uteslutande härledda rättigheter , vilket förstärker deras ekonomiska beroende .
Med tanke på de förändrade ekonomiska och sociala förhållandena bör en av partnern oberoende , individualiserad social trygghet eftersträvas , som garanterar en varaktig trygghet .
Men arbete måste , med alla nödvändiga avgifter , fortfarande också vara lönsamt !
En reform av den sociala tryggheten måste omfatta främjande och försäkringsrättsligt erkännande av tider för barnuppfostran respektive vård av hjälpbehövande familjemedlemmar .
Det alltmer ökande antalet äldre kvinnor som lever i armod är förskräckande .
De kunde genom sin insats för familjen inte prestera någon avgift till det sociala trygghetssystemet ; men även dessa kvinnor måste vara försäkrade .
Ett högvärdigt hälsovårdssystem måste garanteras oavsett den enskildes ekonomiska prestationsförmåga .
Fortfarande är medlemsstaterna principiellt ansvariga för utformningen och finansieringen av sina sociala trygghetssystem .
Men samarbetet inom EU genom expertgrupperna , där naturligtvis kvinnor måste vara rimligt företrädda , kan på lång sikt bidra till en harmonisering av de sociala trygghetssystemen .
Herr talman !
Jag skulle vilja gratulera föredraganden , Andersson , till betänkandet om moderniseringen av den sociala tryggheten som det nu lagts fram .
Som samordnare för Europeiska folkpartiet i utskottet för sysselsättning och socialfrågor är jag mycket glad åt den uppnådda kompromissen som Andersson arbetat så hårt för .
Jag är också mycket glad åt att han fortsatt på ett betänkande jag själv som föredragande skrev i det förra parlamentet och dragen i det här betänkandet är till viss del även samma drag som i det gamla betänkandet .
Syftet med det meddelande från kommissionen i juni 1999 som ligger till grund för Anderssonbetänkandet , är att fördjupa samarbetet mellan medlemsstaterna och EU inom området social trygghet .
Viktiga delmål i detta är : främja sysselsättningen , se till att arbetet ger en fast inkomst .
För det andra , säkerställa pensionssystemen och göra dem betalbara .
För det tredje , främja den sociala integreringen .
För det fjärde , garantera ett betalbart hälsoskydd på hög nivå .
Vid alla dessa målsättningar måste könsrelaterade aspekter spela en viktig roll .
Jag tycker att kommissionen bör lyckönskas till det här meddelandet .
De här fyra punkterna är nämligen mycket viktiga punkter för en hel del medborgare i Europeiska unionen , kanske till och med de viktigaste punkter man funderar över .
Kommissionens meddelande är en viktig strategisk handling för förverkligande av den europeiska sociala konvergensen .
Den makroekonomiska politiken , sysselsättningspolitiken och socialpolitiken påverkas av varandra och måste därför bättre kopplas ihop med varandra .
Kommissionen har insett det sammanhanget .
Meningen är att det åstadkoms en integrerad social strategi som naturligtvis har allt att göra med en bra makroekonomisk strategi och med en bra sysselsättningsstrategi .
De sakerna går inte att skilja från varandra .
Det är endast märkvärdigt att det här förslaget hittills egentligen inte varit en del av en strategi och därför är kommissionens meddelande till viss del ett genombrott .
Något som också är ovanligt glädjande är att rådet nu verkar acceptera det genombrottet och även vill ta upp det i Lissabon .
Vi får naturligtvis inte heller ha för högt uppskruvade förväntningar .
Det är början på en process .
Det är inte slutet på en process .
En del personer har sagt : om vi inte frågar för litet så blir det inte för litet sagt .
Det är dock mycket viktigt att processen kommer igång .
Det rör sig om mycket speciella saker men systemen inom Europeiska unionen är ganska olika .
Utmaningarna är olika .
Arbetslöshetssiffrorna är olika och därför är det mycket viktigt att i det avseendet börja blygsamt men ändå gå vidare ordentligt .
På det sättet kan vi klara en del riktigt stora utmaningar .
I min grupp anser den allra största majoriteten att något sådant måste ske .
Det lustiga med Anderssonbetänkandet är att det inte går in så mycket på diverse detaljer om hur det borde se ut , i det avseendet är det inte ett luftslottsbetänkande .
Det är ett betänkande som försöker visa vägen .
Här och där finns det visserligen några punkter där jag undrar om vi inte är litet för specifika .
Jag tror att en del kolleger kommer att ta upp det igen .
Det hindrar dock inte att det viktiga i betänkandet är att vi utvecklar en strategi , att det finns en rimlig chans att det kan vara ett viktigt bidrag i Lissabon .
Jag tror att om det skulle antas i Lissabon som det ser ut nu så skulle Lissabon bli en stor framgång .
Om det inte antas så säger man i Lissabon egentligen inte så mycket mer än vad som tidigare redan sagts .
I det avseendet är det här betänkandet visserligen bara en del , men kanske den allra viktigaste delen av Lissabonmötet eftersom det verkligen är nytt , medan många andra saker endast är gammalt material i en ny snygg förpackning .
Till sist vill jag hjärtligt tacka föredraganden och utskottet för det här betänkandet .
Jag hoppas att Europa på området social trygghet går ett steg längre med iakttagande av subsidiariteten , för utan den går det inte .
Fru kommissionär , bästa kolleger !
Låt mig , precis som min kollega Bartho Pronk , tacka kommissionen för det här meddelandet och framför allt också gratulera vår föredragande till hans arbete med det här betänkandet .
Det är inte för att det här betänkandet inte längre är kontroversiellt här i parlamentet som det inte skulle vara väldigt viktigt .
Jag har varit med om andra tider då sådana diskussioner om social trygghet egentligen var svåra här i parlamentet .
Diskussionen kommer också alldeles vid rätt tillfälle - Pronk sade det också alldeles nyss - nämligen under förberedandet av toppmötet i Lissabon , där man skall begrunda frågan hur vi via informationssamhället kan ta upp ekonomisk tillväxt , sysselsättning och socialt sammanhang på dagordningen i Europa .
Det är självklart att den sociala tryggheten för min partigrupp är en viktig del av det sociala sammanhanget och därför också måste tas upp på dagordningen i Lissabon .
Min grupp är glad att rådet ( sociala frågor ) redan förra året gav klartecken för en bättre samarbetsstrategi och att en grupp högre tjänstemän förresten redan fått i uppdrag att i juni 2000 lägga fram en första rapport till rådet .
Vi skulle dock som parlament , och framför allt som socialdemokratisk grupp , vilja att Lissabon går ett steg längre .
Det är mycket viktigt att Europaparlamentet i det här betänkandet från vår kollega yrkar för en äkta europeisk strategi med social konvergens , i linje med den så kallade Luxemburgstrategin för sysselsättning , alltså med gemensamma målsättningar , med riktlinjer , nationella handlingsplaner och utvärdering av prestationer .
Vi tycker att den vägen är ambitiös men ändå genomförbar .
Det är naturligtvis självklart att en harmonisering av den sociala tryggheten på europeisk nivå inte är lätt att genomföra .
Systemen för finansiering och organisation är alldeles för olika och det är också ett viktigt skäl till att den sociala tryggheten knappt nått upp på den europeiska dagordningen och att även scenarior som till exempel Danny Peters trettonde medlemsstat eller den europeiska sociala ormen egentligen knappt kommit någonstans .
Den här nya vägen är dock mycket intressant .
Sysselsättningsstrategin har bevisat att den kan fungera och social konvergens behövs också , för våra sociala trygghetssystem står inför samma utmaningar och i EMU-eran riskerar annars alla sociala trygghetssystem att bli en del av den sociala konkurrensen .
Jag vill dock tydligt säga en sak för min grupps räkning : sociala konvergensstrategier får inte bli ett alternativ för social lagstiftning .
De får endast fungera som mycket nyttiga komplement till det vi utarbetar och det vi förväntar från kommissionen med avseende på social lagstiftning .
Jag tror också att det är bra om Europaparlamentet dessutom försöker övertyga rådet att redan i Lissabon konkretisera den samordnade strategin och redan i början av år 2001 inleda ett årligt förfarande för att tvinga tillbaka fattigdomen .
Jag är glad att Europaparlamentet stöder den här idén från min grupp och vi hoppas , fru kommissionär , att vi också kan få ert stöd .
Till sist yrkar vi för att Europaparlamentet och arbetsmarknadens parter och de icke-statliga organisationerna blir nära involverade i den här processen .
Det är endast en bred och demokratisk stödyta som kan ge garantier för att den här strategin lyckas och vi hoppas därför på ert stöd .
Herr talman !
De fyra huvudmål som EU-ländernas regeringar anslöt sig till i november förra året och som nämnts tidigare här i dag , dvs. att man skall se till att det skall löna sig att arbeta och få en fast inkomst , att man skall säkra pensionerna och göra pensionssystemen hållbara , att man skall främja social integration och att man skall se till att få en hållbar sjuk- och hälsovård av hög kvalitet , det är fyra mål som är så brett formulerade att alla bör kunna stödja dem .
Och att låta en grupp höga tjänstemän ha rollen som knutpunkt vid utbyte av erfarenheter för samordning och utvärdering av utvecklingen i social- och arbetsmarknadspolitiken - det kan vi allihop bara bli klokare av .
Kommissionens meddelande som vi diskuterar i dag och som utgjorde grund till rådets beslut i november , är en välbalanserad redogörelse för hur vi kan få en mer kvalificerad debatt , hur vi kan få mer kunskap om de utmaningar som medlemsstaterna står inför på socialpolitikens område under de kommande åren , i och med åldrande befolkning och effekterna av utvidgningen .
Redan i dag har vi stora sociala problem och stora sociala utgifter som belastar de offentliga budgetarna , vilket är ett problem för många medlemsstater .
Sker det ingen reformering riskerar vi att urholka den ekonomiska grunden för socialpolitiken , och en stark och konkurrenskraftig ekonomi är ju den säkraste grunden för en god social trygghet .
Så det är klokt att sätta dessa frågor på dagordningen .
I debatten om samordning av socialpolitiken i EU använder vi ofta uttrycket social konvergens .
Begreppet social konvergens kan vi som liberala ställa upp på när det handlar om att vi i EU fastställer gemensamma , breda målsättningar som länderna försöker uppfylla genom den nationella socialpolitiken .
Det handlar alltså inte om harmonisering , utan om ett gemensamt mål .
Det är ju ett faktum att EU-länderna använder olika sätt att organisera sin socialpolitik .
Vi har olika traditioner , det finns kulturskillnader , och trots många likheter finns det också stora skillnader i de sociala problemens karaktär och i deras omfattning från land till land .
Därför är det viktigt att betona att socialpolitiken är en nationell angelägenhet .
Den nationella politiken är naturligtvis styrd av en rad gemensamma ramar som gäller de sociala minimirättigheterna , som regleras i fördraget , rörande hänsynen att vi skall samordna ekonomierna och det ekonomiska samarbetet .
Det skall alltså vara en samordning och ett samarbete .
Men konvergensen gäller målen , inte medlen .
Jag vill också gärna tacka föredraganden , Jan Andersson , för betänkandet och för hans mycket konstruktiva insats för att försöka sammanjämka olika ståndpunkter och säkerställa ett stöd till sitt betänkande .
Jag kan stödja betänkandet , men det finns enskilda punkter som inte är helt i min smak .
Jag stöder inte kravet på att kommissionen skall ingripa vid s.k. orättvis konkurrens mellan social- och skattesystem , om ett sådant ingrepp skall användas för att hindra nytänkande , utveckling och effektivisering av våra sociala system , eller användas för att hindra en sänkning av det alltför höga skattetrycket i många EU-länder .
Jag är skeptisk rörande den detaljreglering som skulle kunna bli resultatet av att kommissionen skall bedöma omfattning och kvalitet i barn- och äldreomsorgen och skeptisk rörande värdet av en gemensam fattigdomsgräns .
Samordning av socialpolitik och dialog är bra , men vi skall inte dra alla över en kam ; det skall finnas utrymme för en mängd olika lösningar .
Herr talman , fru kommissionär !
I samband med den strategi för modernisering av den sociala tryggheten som förklarats här , vill jag ändå ta upp några punkter , några positiva och några frågetecken .
Jag är positiv till att det här ärendet sakta men säkert satts i rörelse .
Det är bra , tycker jag .
Det verkar vara nyttigt .
Jag kan också vara positiv till de stora dragen i meddelandet , det strategiska handlingssättet .
Vi hoppas därför också att de fyra målsättningar som nämns här också kan uppnås på ett rimligt sätt .
Vi vill också betona vikten av hur det hanteras , å ena sidan processen à la Luxemburg , riktlinjer , men vi tror också att det är viktigt att , som Van Lancker redan sagt , det ställs upp riktlinjer för till exempel atypiskt arbete , enmansföretag , och så vidare .
Vi urskiljer dock två problem som vi måste försöka hitta lösningar för .
Det första är att det talas om att anpassa den sociala tryggheten nedåt , när vi hoppas att det talas om konvergens på samma nivå .
Jag skall ge några exempel från en undersökning som den nederländska fackrörelsen nyligen genomförde angående reformerna i Europeiska unionen med avseende på den sociala tryggheten .
Där visar det sig att anpassningar går att hitta överallt .
Många av de anpassningarna , majoriteten av dem till och med , visar sig dock vara anpassningar nedåt , resten är förbättringar .
Majoriteten av de anpassningarna är inriktade på pensioner , elva inskränkningar och två förbättringar .
När det gäller arbetslöshetsersättningen finner vi sex inskränkningar och fem förbättringar .
Skälen till anpassningarna är till exempel förbättring av sysselsättningen , minskning av utgifterna för den sociala tryggheten men även politisk konkurrens och EMU-kriterierna .
Den politiska konkurrensen finner vi främst i de nordliga länderna .
Den mesta stabiliteten och till och med förbättring av den sociala tryggheten ser vi i de sydliga länderna .
Sammantaget ser vi också en begränsad roll för arbetsmarknadens parter i hela den här processen .
Det är inte glädjande och betyder att konvergensstrategin måste inriktas på de bästa handlingssätten .
Cappuccino , för att uttrycka det så , är inte alltid välgörande för oss .
Herr talman !
Jag kommer från samma land och samma region som föredraganden Andersson .
I min valkrets finns det en djup skepsis mot kommissionens styrnings- och kontrollförsök .
Om Anderssons väljare visste att han föreslår att socialpolitiken i hela Europa skall samordnas , att skatterna skall harmonieras och att välfärdssystemet skall inordnas under EMU-processen , skulle de protestera högt och tydligt .
Jag är säker på att de flesta skulle rösta på ett annat parti nästa gång .
Visserligen har Anderssons betänkande många bra konkreta förslag , som jag kan stödja helt och hållet .
Jag är dock kritisk till det helhetsperspektiv för social trygghet , som präglar både kommissionens meddelande och Anderssons betänkande .
De tycks tro att det är kommissionen som är motor , centrum och drivkraft i förändringsprocessen i Europa .
Precis som Prodi i förmiddags beskrev sig själv som en person som bär all världens ansvar på sina axlar , så möter vi här ett uppifrån-perspektiv på de sociala frågorna .
Man talar om konvergens och harmonisering med detta uppifrån-perspektiv .
Man försöker till och med få oss att tro att social integration kan tänkas vara en gemensam alleuropeisk process .
Verkligheten är helt annorlunda .
Ett socialt integrerat Europa är en avlägsen utopi , som inte ens en allsmäktig kommission kan förverkliga .
Man har tagit stora steg mot ekonomisk integration .
Man är i färd med att skapa en politisk integration .
Men social integration är ett helt annat slags process , som förutsätter kulturell gemenskap och direktkommunikation mellan människor .
Idén om det sociala Europa är en skrivbordsprodukt , som är långt från verklighetens värld .
Socialpolitiken är i huvudsak en nationell process .
I mitt hemland har vi lärt oss att stora delar av den sociala tryggheten måste skapas lokalt inom kommunernas ram .
Decentralisering och närhet är viktiga för kvalitet och effektivitet inom vård , skola och sociala tjänster .
Kommunerna har ansvaret för nästan all produktion av välfärdstjänster .
Den kommunala demokratin är ramen för social trygghet .
När vi nu har fått en ekonomisk samordning , tror jag visserligen att det behövs en växande grad av samordning av även socialpolitiken på europeiskt plan .
En europeisk strategi för samordning måste bygga på lokala initiativ , på mångfald .
Den måste respektera närhetsprincipen och vara demokratiskt förankrad .
Jag tillhör ett parti som en gång trodde på central styrning , femårsplaner och långtgående konvergenskrav .
Vi tog gruvligt fel och historien tvingade oss till självkritik , omtänkande och andra föreställningar om demokrati .
Jag tror inte att huvudansvaret kan vila på Prodi och hans kommission .
Jag är övertygad om att det måste bäras av de människor som är direkt berörda av de sociala problemen .
Herr talman !
Jag skulle i min tur vilja gratulera både kommissionen och föredraganden .
Kommissionen eftersom ett nytt steg tagits i konvergensen mot social trygghet och föredraganden för det goda betänkande han utarbetat .
Europeiska unionens politik omfattar förutom en ekonomisk politik och en sysselsättningspolitik även en socialpolitik .
Hittills har den varit begränsad , både när det gäller utformning och medel .
Under inflytande av den fria rörligheten för arbetstagare , av den inre marknaden och av euron så integreras dock även arbetsmarknaderna .
Det har utan tvekan konsekvenser för den sociala tryggheten som i stor utsträckning är bunden till arbete .
Gränsarbetare , utstationerade arbetstagare , utflyttade arbetstagare men även arbetssökande , praktikanter och studenter ser sig förhindrade att utöva rätten till fri rörlighet och det till följd av bristen på samordning och avsaknaden av konvergens i den sociala tryggheten .
Samma fenomen förekommer förresten också inom skatteområdet .
För att bekämpa både konkurrensstörningar och dumpning så har kommissionen så vitt jag kan se utvecklat ett tillvägagångssätt som balanserar mitt emellan å ena sidan harmonisering och å den andra sidan icke-inblandning .
Å ena sidan använder man bindande och framtvingbara regler för lika löner eller för kompletterande pensioner och å andra sidan använder man program för att ge stimulans med avseende på icke-diskriminering eller social utslagning .
På grundval av en serie rekommendationer , rapporter och meddelanden har kommissionen tagit ett extra steg i riktning mot konvergensen , nämligen genom att å ena sidan sätta upp målsättningar och å den andra inrätta en arbetsgrupp med topptjänstemän .
Båda förslagen har redan accepterats av rådet och det gäller alltså att stödja det tillvägagångssättet för att på sikt , med sakkunskap , kunna bedöma om och i vilken utsträckning och på vilket sätt den sociala tryggheten i Europeiska unionen måste omorganiseras .
Utvidgning , globalisering , åldersökning , individualisering och familjeförändringar gör en sådan omorganisering oundviklig .
Att förneka dessa förändringar är egentligen detsamma som att ge upp den sociala tryggheten .
Till EU-skeptiker och nationalister säger jag att en social trygghet som endast gäller innanför medlemsstatens gränser inte är social och inte ger något skydd .
En nedrustning på grund av konkurrens till den sociala tryggheten skadar nämligen samtidigt den sociala tryggheten som produktiv faktor .
Mindre social trygghet betyder också mindre köpkraft , färre friska arbetstagare och färre lyckliga arbetstagare .
Till supereuropéerna säger jag att en europeisk social trygghet inte är genomförbar och inte heller önskvärd .
Skillnaderna mellan medlemsstaterna är alldeles för stora , både när det gäller faciliteter , berättigande , inkomster och utgifter , osv .
Ett jämställande är alltså omöjligt att genomföra .
Den väg som kommissionen följer är faktiskt självklar .
Fördelarna är tydlighet , insamling av uppgifter , utbyte av erfarenheter för att sedan komma överens och ställa upp indikatorer för jämförelse och ge rekommendationer .
Jag ställer mig bakom den uppfattningen .
Jag stöder kommissionen och jag hoppas att Lissabon i det avseendet tar ytterligare ett steg framåt .
Jag vill tacka föredraganden för det berikande bidraget till kommissionens initiativ .
Trots viss skepticism hos några så är vi överens om att vi måste ha en fast strategi för att förnya det sociala skyddet .
Åttio- och nittiotalets debatter visar vikten av social transferering .
Mer än 50 procent av unionens medborgare mottar förmåner som inte härrör från pensioner .
Danmark och Nederländerna är positiva exempel på hur vi alla måste anstränga oss för att få sammanhållning .
Mer än 60 procent av de medborgare som befinner sig i farozonen har i de här länderna tagit sig ur fattigdom .
I länderna i söder är det däremot bara mellan 7 och 15 procent som klarar av det .
Detta genererar social orättvisor och den redan nämnda konkurrensen .
Konvergenskriterierna fick oss att dra ned på de offentliga utgifterna , vilket ledde till en anti-europeisk stämning .
Sanningen är att höga skyddsnivåer går hand i hand med högre produktivitet .
En konvergensstrategi för den sociala politiken , som åsyftas i betänkandet , kan också vara fördelaktigt för medborgarna och för den inre marknaden .
Alla system stöter på nya problem , vilka identifieras i betänkandet .
Den demografiska frågan är central , men nya arbetsformer , rörligheten inom unionen , kortare aktivt liv ( dagens ungdom kommer senare till arbetsmarknaden och man har föregripet reformen om lagliga 65 år till faktiska 57 / 59 år på grund av industriella omstruktureringar ) är också viktiga frågor .
Att fattigdomen är ett ihållande fenomen blir man mer och mer medveten om , särskilt för kvinnorna i reformen , tack vare låga löner och otillräckliga bidrag .
Utmaningar som dessa måste få ett snabbt svar .
Det portugisiska ordförandeskapets initiativ är mycket välkommet : att inrätta en grupp på hög nivå , den nivå vi vill att lagstiftande åtgärder skall förberedas och utarbetas på .
Problemet skall inte bara skjutas upp eller ställas en simpel diagnos på .
Vi behöver gemensamma , temporärt realistiska mål vid horisonten .
Herr talman !
Anderssons betänkande innehåller mycket av intresse .
Tyvärr är dock det mest intressanta att betänkandet , som skall antas behandla en samlad strategi för en modernisering av socialpolitiken , i stället föreslår en utbyggnad av traditionell socialpolitik och mer överstatlighet på det sociala området .
Socialpolitiken måste förnyas för att arbetslösheten i medlemsstaterna skall kunna minskas .
Även om socialisterna , när det numera finns så många socialdemokratiska regeringar , talar mycket mindre om arbetslösheten än tidigare , är denna arbetslöshet förfärande hög .
Detta trots en internationell högkonjunktur .
Något måste göras för att arbetslösheten inte skall förvandla den så kallade europeiska modellen till en parodi .
Socialpolitiken måste underlätta sysselsättning , skapa incitament till ökad sysselsättning både hos arbetsgivare och arbetstagare .
I Anderssons betänkande krävs social konvergens , det vill säga att systemen alltmer skall likriktas inom och genom EU .
EU skall anta , som det heter , verkliga konvergenskriterier , som är bindande och effektiva .
Andersson vill också ha en effektiv och ambitiös skattesamordning , det vill säga överstatlighet på skatteområdet .
EU skall också , på grundval av en enhetlig definition av fattigdomsgränser , lägga fram rekommendationer om vad som kallas godtagbart minimiuppehälle i medlemsstaterna .
EU skall arbeta fram riktlinjer för kvaliteten i de arbetstillfällen som skapas , vad nu det kan betyda .
Inte kommer arbetslösheten att kunna minskas med alla dessa ytterligare regleringar och ingrepp .
De strukturella problem , som gör arbetslösheten högre i Europa än i Förenta staterna , kommer att bli ännu större .
Det behövs ingen överstatlighet på det här området .
Medlemsstaterna kan utforma sina egna system på det sociala området , var och en inom ramen för sina ekonomiska resurser och politiska preferenser .
Detta är alldeles särskilt viktigt för att inte skapa onödiga problem inför utvidgningen av EU .
Andersson menar att de fattiga östländerna skall påminnas om att den sociala konvergensen skall omfatta även dem .
Det är dock uppenbart att dessa länder , utarmade inom ett kommunistiskt ekonomiskt system , inte kan hålla sig med en socialpolitik som till exempel Sveriges .
Minimiregler och fattigdomsgränser blir antingen meningslösa för de nuvarande medlemsstaterna eller orimliga för fattiga kandidatländer .
Herr talman !
Jag vill liksom övriga också gratulera Andersson till hans betänkande .
Han har utfört mycket arbete för parlamentets räkning för att ta fram en bred samsyn om vad som definitionsmässigt är en kinkig fråga inte bara i detta parlament utan i praktiskt taget varje medlemsstat .
Jag är också positiv till kommissionens meddelande .
Den lät vänta på sig men väl värd att vänta på .
Det kan bli ett landmärke för utvecklingen av ett socialt Europa , under förutsättning av vi menar allvar och inte tillåter enskilda medlemsstater att rygga för de åtgärder som måste vidtas för att genomföra det .
Vi kan och måste ta den unika europeiska samhällsmodell vi har och omforma den för att passa in i 2000-talet , ett århundrade där en snabb globalisering sker .
Jag är rädd för att de förslag som lagts fram av Herman Schmid inte tar upp den globaliseringen i världen .
För att lyckas måste vi se till att vår ekonomiska politik , vår sysselsättningspolitik och vår politik för social trygghet i dess vidaste mening integreras och av vi hanterar dem som en helhet .
Vi måste se till att våra Ekofin-ministrar och våra arbetsmarknadsministrar tillstår att socialministrar kan medverka i arbetet med att upprätta ett samhälle i Europa som är kreativt , initiativrikt och som skall höja alla våra medborgares livskvalitet .
Detta är inte längre fråga om ett val för oss .
Det är en tvingande nödvändighet .
Europas medborgare kommer inte att nöja sig med mindre än en livskvalitet som gagnar dem som människor .
Vi vill inte ha den amerikanska modellen - en modell som har misslyckats att skapa den sysselsättningsnivå som krävs för att ge en anständig livskvalitet .
Vad den har resulterat i är en dramatisk ökning av fattiga arbetstagare i Förenta staterna .
Det är inte vad vi vill göra i Europa .
Vi har en tradition av solidaritet i Europa och vi har erfarenhet av ett bättre sätt att göra saker .
Men vi måste få tag i verktygen för att göra detta .
Jag yrkar därför på att vi inte bara inrättar den arbetsgrupp på hög nivå som kommissionen föreslagit utan också går vidare och genomför en typ av Luxemburgprocess så att vi får en integrerad strategi för denna fråga om social trygghet .
Herr talman , ärade kommissionär !
Det här är ett av de sociala områden som Europeiska unionen borde uppmärksamma betydligt bättre .
Sanningen är att den makroekonomiska politiken , stabilitetspakten och de nominella konvergenskriterierna har bromsat förnyelsen av det sociala skydd som bidrar till bättre livskvalitet hos befolkningen , främst genom starkt höjda pensioner och andra reformer , särskilt minimipensionerna , och kampen mot socialt utanförskap .
Detta är särskilt allvarligt i länder som Portugal , där pensioner och minimireformer knappt uppgår till hälften av den nationella minimilönen , vilken i sin tur är den lägsta i hela Europeiska unionen .
Förstår inte kommissionen vikten av att ändra på den makroekonomiska politiken för att skapa kvalitativ sysselsättning med rättigheter , grundläggande för att bevara och modernisera ett starkt system för det offentliga sociala skyddet , så tvivlar vi starkt på deras ståndpunkt .
Trots att man i Andersonbetänkandet tog upp en del positiva förslag , några av dem som vi hade lagt fram , kvarstår delar av den grund vi kritiserade i kommissionens förslag och den oro vi känner inför strategin för en reformering av det sociala skyddet .
Herr talman !
I mitt tidigare arbetsliv skötte jag två produktionsföretag , ett i Förenade kungariket och ett i Nederländerna .
När företaget i Förenade kungariket växte investerade vi i mer personal , när det holländska företaget växte investerade vi i fler maskiner .
Det enkla skälet till detta var att de sociala kostnaderna i Nederländerna var alltför höga vid en jämförelse .
Jag är positiv till social trygghet , jag är positiv till kommissionens ursprungliga dokument men jag önskar inte se människor förlora jobben på grund av att socialförsäkringskostnaderna blir orealistiskt höga .
Det var därför jag i utskottet föreslog någon form av utvärdering av effekten på företag så att hänsyn kunde tas till kostnader och risker för sysselsättningen och EPP-DE gruppen stödde detta ändringsförslag .
Men jag måste konstatera att andra grupper , ledda av PSE-gruppen och min landsman , Stephen Hughes , röstade emot detta .
Jag håller med om att Anderssons betänkande är mycket välmenande och jag högaktar honom för det arbete han har gjort men enligt min mening skulle det sätt som social konvergens definieras och stöds i betänkandet innebära att man driver upp samhällskostnaderna till högre nivåer i hela EU .
Det skulle leda till att flera jobb hamnar i riskzonen och även riskera denna kammares trovärdighet genom att spegla hur fjärran vi befinner oss från den verkliga världen .
Jag uppmanar därför denna kammare att avslå hela betänkandet och låta det ursprungliga förslaget från kommissionen , som var mycket väl avvägt , fortfarande gälla utan ändring .
Herr talman , vi kan inte rösta för detta betänkande .
Europeiska unionen bör sätta det sociala i centrum för uppbyggnaden .
Det är de sociala rättigheterna som borde styra ekonomiska val och inte tvärtom .
Därför när det gäller det sociala trygghetssystemet är vi emot införandet av mekanismer som kopieras på Luxemburgprocessen och går emot denna tanke : stora ekonomiska riktlinjer , sedan konvergenskriterier och slutligen det sociala som behandlas som en restvara .
Europeiska unionen borde proklamera en allmän princip : de sociala rättigheter som uppnåtts i staterna kan inte minskas .
Varje insats av gemenskapen borde syfta till att komplettera och sedan harmonisera uppifrån de befintliga garantierna .
För att stärka finansieringen av de sociala trygghetssystemen behövs det en allmän löneökningspolitik och införandet av ett lagenligt lägsta lönetak i alla medlemsstater .
För att bekämpa fattigdom är rätt till inkomst och rätt till sysselsättning oskiljaktiga .
För att till slut undvika att hälsovården behandlas som en vara bör Europeiska unionen uttala sig klart och tydligt mot pensionsfonder och sätta sig upp emot att privata försäkringsbolag har tillträde till hälsovårdssystemet .
Avslutningsvis tror jag verkligen att ett socialt Europa inte kan nöja sig med uttalanden och fromma önskningar .
Läget är alltför tragiskt för miljoner människor .
Herr talman , fru kommissionär , ärade ledamöter !
Målsättningen att skapa en samordnad strategi för att modernisera den sociala tryggheten inom Europeiska unionen är helt klart någonting positivt .
Det var också positivt att man , i och med toppmötet i Luxemburg , drog igång den europeiska strategin för samordning av sysselsättnings- och arbetsmarknadspolitiken .
Arbetsmarknad och social trygghet är egentligen två sidor av samma sak , och kräver synkroniserad politik och reglering .
Om arbetsmarknaden fungerar vad sysselsättningsnivåer , flexibilitet och löneeffektivitet beträffar , fungerar också välfärdsstaten och den sociala tryggheten och vice versa .
Fram till helt nyligen fastställde Europas länder internt , på ett så att säga självförvaltande sätt , reglerna för hur dessa två marknader skulle fungera och finansieras .
Budget- och växelkurspolitiken sörjde för intern och extern balans .
I och med Maastricht och den gemensamma valutan blev budgetpolitiken starkt kringskuren och man kan inte längre ta till devalvering i jakten på förlorad konkurrenskraft .
De strukturella och konjunkturmässiga klyftorna mellan länderna kan därför inte överbryggas med hjälp av underskott och växelkurser .
Eftersom läget är sådant är det bara arbetsmarknaden och välfärden som kan stå för en flexibilitet för att avhjälpa både de strukturella och de konjunkturberoende obalanserna , de så kallade asymmetriska esogena chockerna , i avsaknad av en full rörlighet för arbetskraft inom unionen och en fördelningspolitik på federal nivå .
Och detta är det paradoxala .
Samordningen av politik och penningmarknad i Europa medför oundvikligen en samordning av spelreglerna för arbetsmarknaden och välfärden , men samtidigt tvingar oss den gemensamma valutan och bristen på arbetskraftsrörlighet och en omfördelande skattepolitik till icke samordning i löne- och välfärdsmässiga termer för att kompensera för olika produktivitetsmarginaler på nationell och regional nivå .
Dessa motstridigheter kommer man inte ur med hyckleri och vackra ord som samordning , benchmarking , modernisering och medlingsförfarande .
Antingen blir Europeiska unionen en riktig federal stat med en riktig fördelningspolitik , en riktig rörlighet för arbetskraften och därmed , först därefter , med gemensamma regler om arbetsmarknad och välfärd , eller också är det bättre att inte bedra eller bedra sig med omöjliga vägar till samordning som låter bra men som i verkligheten skadar framför allt de svagaste .
Och det vore bra om alla vore medvetna om detta .
Herr talman !
I motsats till mina kolleger i dagens debatt är jag böjd att rösta för Anderssons betänkande , bl.a. därför att jag ser mycket tydliga skillnader jämfört med kommissionens meddelanden .
I synnerhet anser jag att detta betänkande - och det vill jag gratulera föredraganden till - försvarar den solidariska ansatsen i den europeiska trygghetsmodellen .
Jag vill framhäva de klara ståndpunkterna mot social dumpning , liksom rätten till social grundtrygghet , målet med den sociala konvergensen och särskilt det som i mycket konkret form , när det gäller kvinnors jämställdhet , har nämnts som mål för socialpolitiken .
Jag ser också de brister som uppstått på grund av en inte tillräckligt konsekvent uppgörelse med den makroekonomiska politiken i Europeiska unionen , som står i vägen för detta solidariska förnyande av den europeiska socialstatsmodellen , men allt som allt ser jag positivt på detta betänkande .
Herr talman !
Jag tar till orda för att påtala och bekräfta behovet av en modernisering av den sociala tryggheten som ett instrument som är mycket mer än ytterligare ett steg mot byggandet av Europa .
Det kommer till uttryck i Anderssons betänkande som jag anser vara alldeles utmärkt .
Europa , Europeiska unionen kommer , även om den ekonomiskt och politiskt sett är stark , att halta , bli försvagad och begränsad , kanske kortlivad , om vi inte har förmåga att stärka den på det sociala området .
Det senare förutsätter , vad jag kan förstå , möjligheter till arbete för dem som kräver detta , men även ett beslutsamt agerande till förmån för de socialt utsatta .
Om man utgår från att alla människor har rätt till en social trygghet och en garanterad minimiinkomst , är det en situation vi inte får glömma bort : situationen för dem som inte är födda i Europeiska unionen .
Låt oss inte glömma att det under 1999 var 717 000 som kom och jämnade ut våra låga födelsetal .
Därför är det helt nödvändigt att den sociala ordningen inbegriper en invandrarpolitik med en social medvetenhet , precis som president Gutierres nyligen sade i Spanien .
Det är viktigt att stor hänsyn tas till situationen för de personer som inför ekonomiska förändringar , sammanslagningar , övertagande , ny teknik , etc. ser sina möjligheter till arbete hotade eller begränsade .
Här krävs en politik med anpassade och förberedande utbildningar till nya arbetstillfällen , för säkrandet av en redan existerande anställning eller för en andra chans , för postmannen ringer alltid på två gånger , för att använda den kända filmens titel .
Jag vill i all anspråkslöshet säga att detta åligger alla europeiska regeringar , såväl på nationell som regional nivå , att se till att han ringer på mer än en gång .
Jag anser , fru kommissionär , att det är kommissionen som bär ansvaret för att initiera och samordna dessa möjligheter .
Herr talman !
Jag skulle vilja gratulera herr Andersson till hans utomordentligt goda arbetsinsats .
Det råder därför ett mycket brett samförstånd , och jag skulle vilja tacka parlamentsledamöterna för deras insatser .
Först vill jag påpeka att de europeiska organen började diskutera de sociala trygghetssystemen redan för ganska många år sedan , och redan 1995 kom den första rapporten med titeln " Den sociala tryggheten i framtiden " .
Det har också kommit betänkanden från Europaparlamentet , från Weiler och Pronk .
I dag behandlar vi Anderssons betänkande .
Jag anser att vi har gjort betydande framsteg , eftersom vi nu talar om en modernisering av de sociala trygghetssystemen .
Den andra punkt jag vill ta upp är att vi måste ta hänsyn till vilken rättslig grund som kan gälla för Europeiska kommissionens verksamhet .
Ni vet mycket väl att fördraget inte innehåller någon rättslig grund för politik på europeisk nivå , däremot finns det en överenskommelse som kom till uttryck också vid det senaste rådsmötet , det finns en överenskommelse om att medlemsstaterna skall inleda ett samarbete , genom samordning och genom erfarenhetsutbyte kring framgångsrika program .
Mitt tredje påpekande gäller följande : betänkandet är koncentrerat till fyra områden ; förvärvsarbete , pensionssystemens hållbarhet , den sociala integrationen och slutligen hälso- och sjukvårdens kvalitet .
På alla dessa områden beaktas kvinnornas situation , eftersom det ­ såsom de kvinnliga parlamentarikerna påpekat ­ inom vart och ett av dessa områden finns speciella problem som gäller kvinnor , och dessa problem bör i många fall lösas genom särskilda politiska insatser .
Nästa punkt gäller de konkreta insatser som vi har gjort .
Som ni vet , har det portugisiska ordförandeskapet redan tillsatt en arbetsgrupp på hög nivå , som kommer att lämna sin första rapport vid toppmötet i juni .
Det portugisiska ordförandeskapet koncentrerar sig på två frågor , långsiktigt hållbara pensionssystem och social integration .
Det är mycket positivt att man föreslagit inrättandet av en motsvarande grupp på parlamentsnivå .
Sedan denna grupp på hög nivå godkänts , kommer vi att kunna gå vidare till nästa steg .
När det gäller de sociala trygghetssystemens roll och kostnaderna för den sociala tryggheten men också den roll som dessa system spelar i konkurrensen mellan medlemsstaterna , skulle jag vilja påpeka att den europeiska politikens strävan är att kombinera konkurrenskraft och social sammanhållning .
Vi måste naturligtvis ta hänsyn till konkurrensaspekten , men när man planerar de sociala trygghetssystemen , måste man se till att den sociala tryggheten blir en viktig faktor för ekonomisk tillväxt och sysselsättning .
Och jag anser att detta klart framgår av innehållet i meddelandet .
Värderade kolleger !
Vårt mål är att vi under nästa år , efter ett enhälligt beslut av rådet , skall kunna åstadkomma samordning , erfarenhetsutbyte , kartläggning av de sociala problemen , en faktabas för att bättre kunna samordna de politiska insatserna .
Såsom många parlamentsledamöter framhållit , tror också jag att vi har tagit ett första , betydelsefullt steg .
Under regeringskonferensen har de socialpolitiska frågorna redan behandlats utifrån ett vidare perspektiv , och jag tror att vi har kommit in i en ny fas , där socialpolitiken i betydande utsträckning kommer att vara en europeisk politik .
Tack , fru Diamantopoulou .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.30 .
 
WIPO-avtalen Nästa punkt på föredragningslistan är rekommendation ( A5-0008 / 2000 ) av Cederschiöld för utskottet för rättsliga frågor och den inre marknaden om förslag till rådets beslut om bemyndigande att på Europeiska gemenskapens vägnar underteckna WIPO-avtalet om upphovsrätt och WIPO-avtalet om utövande konstnärer och ljudupptagningar ( KOM ( 1998 ) 249 - C5-0222 / 1999 - 1998 / 0141 ( AVC ) ) . .
Herr talman !
Vi tar nu ställning till en viktig fråga , ett internationellt avtal , en fråga som kan komma att påverka välståndsutvecklingen i många medlemsstater .
I mitt hemland , Sverige , berörs en av de största exportbranscherna .
Musik och ljudupptagningar är områden som berörs .
Det handlar om konstnärers rätt till upphovsrätt , till skydd för sina konstnärliga produkter .
Det handlar om WCT ( World Copyright Treaty ) och WPPT ( World Perfomance and Phonograms Treaty ) .
Utan immaterialrättsligt skydd hämmas de ekonomiska incitamenten och skaparkraften .
Förfalskningar är big business .
Man räknar med att man bara i Europa går miste om inkomster på 4,5 miljarder euro på grund av piratkopiering .
Problemet berör många arbetstillfällen i underhållningsbranschen .
Detta är ett historiskt avtal , eftersom EU är fördragsslutande part .
Så är fallet trots att inte EU , utan endast medlemsstaterna , är med i organisationen .
Det finns en särskild klausul , som kräver parlamentets samtycke i två fall .
Vad gäller detta avtal är båda dessa villkor uppfyllda .
Det skapas en ny institution , en församling som fortsättningsvis skall följa upp avtalet och dess konsekvenser .
Dessutom berör avtalet frågor , som behandlas i enlighet med medbeslutandeförfarandet .
Parlamentet måste således ge sitt samtycke , eftersom det berör dess kompetens .
Framtiden kommer att utvisa om det är riktigt att genom denna nya parlamentariska församlingen skära ner kommissionens kompetens i dessa frågor .
Parlamentet kan i varje fall för närvarande inte göra något åt saken .
Avtalet kompletterar Bern-konventionen , när det gäller litterära verk .
Ett internationellt rättsligt skydd skapas för spridning , försäljning , uthyrning , offentlig återgivning och tillhandahållande .
Dessutom skapas skydd för programvaror och databaser .
Problem föreligger när det gäller begreppet " upphovsman " .
Det är till exempel inte definierat .
En annan fråga , som utgör ett visst problem , är frågan om mellanlagringar .
Den är inte heller löst .
Den behandlas genom en generalklausul , som inte har någon definition .
Om man inte gör några preciseringar i denna typ av frågor , kan det leda till att de hanteras olika runt om i världen , utan enhetlighet .
Detta skulle inte vara bra .
Frågan om skiljedomsprövning återstår också att lösa .
Parlamentet kan inte ändra dessa enskildheter .
Vi kan bara säga ja eller nej till avtalet , som det föreligger - ja eller nej till ett avtal med brister .
Både jag , som föredragande , och utskottet tycker att vi bör säga ja .
Vi har här ett avtal som trots sina brister innebär ett betydande steg framåt för upphovsrätten .
Vi har ju länge diskuterat om parlamentet och om EU skall ha kompetens när det gäller patentfrågorna i immaterialrätten .
Jag tycker det .
Det finns dock ännu ingen gemenskapslagstiftning på området patenträtt och mönsterskydd , men det behövs .
Ett europapatent är på väg , vilket är bra .
Nu tar unionen och medlemsstaterna tillsammans de första stegen på det immaterialrättsliga området .
Det är bra för oss om vi har kraften att göra det , trots att vi inte är helt nöjda .
Vi kan därigenom fungera som en förebild för kandidatländerna .
Vi har ett direkt ekonomiskt intresse av att dessa frågor regleras före utvidgningen .
Jag vill tacka kommissionen för insatserna på området och för samarbetet med kommissionens tjänstemän , som har varit alldeles utmärkt .
Till sist vill jag tacka även kammaren för att man varit vänlig och åhört dessa ord vid denna sena timme .
Herr talman !
Också jag skulle vilja gratulera föredraganden Cederschiöld till en mycket betydelsefull arbetsinsats .
Hon har tydligt klargjort de problem som uppstår genom godkännandet av WIPO-avtalet .
Godkännandet av avtalsvillkoren är otvivelaktigt en historisk händelse , eftersom Europeiska unionen för första gången medverkar som avtalsslutande part i ett internationellt avtal på det immaterialrättsliga området .
Vägen dit har verkligen varit lång , främst på grund av den juridiska frågan om i vilken mån gemenskapen skulle kunna anses ha fullständig behörighet i fråga om immaterialrätt .
Problemet har nu lösts .
I dag uppmanas vi att ge vårt samtycke till vad som egentligen är två avtal : avtalet om immaterialrätt och avtalet om tolkningar , framföranden och ljudupptagningar .
Det första avtalet förefaller på ett effektivt sätt uppfylla de krav som ständigt framförts av upphovsmän till konstnärliga och litterära verk , samtidigt som det ger ett skydd i fråga om spridning , uthyrning och offentligt återgivande av konstnärers och författares verk .
I fråga om det andra avtalet , som gäller framföranden och ljudupptagningar , bör det framhållas att det är första gången som ett internationellt avtal , undertecknat även av gemenskapen , erkänner utövande konstnärers exklusiva rätt till kopiering , spridning och uthyrning av sina verk till allmänheten samt rätten till skälig ersättning för radioutsändningar .
I fråga om kopieringsrätten innebär avtalet ett betydande framsteg .
Kommissionen påpekar att det i avtalstexterna inte finns några specialbestämmelser som täcker alla frågor som uppstår genom den tekniska utvecklingen .
Ändå kan man hävda att de utövande konstnärerna genom avtalen får ett bättre rättsligt skydd än de tidigare haft med stöd av Romfördraget eller av gemenskapens olika direktiv .
Den slutsats jag drar av artikel 7 i avtalet är att kopieringsskyddet inte bara gäller de framföranden som finns på ljudupptagningar och som framförs av de utövande konstnärerna själva , utan alla typer av kopiering , delvis eller fullständig , lång- eller kortvarig , och alla andra typer av produktioner .
Jag vill emellertid också lyfta fram ett antal punkter som bör uppmärksammas vid kommande WIPO-överläggningar eller andra diplomatiska överläggningar .
Det gäller först rätten till spridning i enlighet med artikel 8 , första stycket .
I nästa stycke i samma artikel ges staterna rätt att återkalla denna rättighet .
Detta är farligt , och det är ett av de mest negativa inslagen i avtalet , eftersom ingenting hindrar staterna att införa specialbestämmelser om upphävande av denna rättighet , vilket skulle få negativa konsekvenser för konstnärerna .
Beträffande rätten till uthyrning tolkar jag artikel 9 så att den exklusiva rätten till uthyrning tillkommer de utövande konstnärerna , om detta föreskrivs i den nationella lagstiftningen , och här anser jag att det finns en skillnad i förhållande till artikel 13 .
Avslutningsvis vill jag säga att dessa avtal öppnar nya perspektiv för upphovsrätten .
Under det tjugoförsta århundradet , kunskapens och den immateriella ekonomins århundrade , kommer immaterialrätten att vara en dominerande ägandeform och i många fall viktigare än det traditionella ägandet .
Vi befinner oss i början av en epok då det kommer att skapas ett nytt rättssystem , i vilket upphovsrätten kommer att vägas mot det offentliga intresset att en bred allmänhet får tillgång till den immateriella egendomen .
Herr talman !
Tack så mycket också till föredraganden !
Jag tror att hon har tagit upp ett par viktiga punkter , som jag också strax kommer att tala om .
Till att börja med diskuterar vi parlamentets godkännande av de nämnda fördragen som hör till WIPO .
Ännu har ingenting trätt i kraft , Europaparlamentets beslut har alltså betydelse denna gång .
EU : s tillträde motsvarar dess önskan att dra till sig all internationell och intern behörighet , men det är oklart var de behörigheter skall ligga som dras bort från den nationella kontrollen .
Ett godkännande kan här alltså bara rekommenderas om Europaparlamentet vid varje vidare utveckling av WIPO-rätten är med från början till slut och har medbeslutanderätt .
Det är inte föreskrivet i Amsterdamfördraget .
Vad säger kommissionen om detta ?
Väsentliga aspekter är fortfarande oklara i förslagen till WIPO-avtalet , det säger även föredraganden .
För att nämna ett exempel : Begreppet " upphovsman " är inte alls definierat i avtalet .
Därigenom skulle rättstvister mellan fördragsparterna vara förprogrammerade .
Här vill jag fråga kommissionen : Vill den gå in med förbundna ögon i detta problem ?
Vill den tvinga på andra avtalsparter sina definitioner av upphovsrätt ?
WIPO : s idé stöder sig också på konceptet om individens rätt .
Det leder t.ex. för urspungsfolket samerna till problem , eftersom de har en annan rättsförståelse , en kollektivrättsförståelse .
Men det är också offentliga intressen som står på spel .
Det är t.ex. oklart om det för offentliga bibliotek i framtiden överhuvud taget fortfarande kommer att vara tillåtet att gratis låna ut böcker , videoband och kassetter .
Härigenom berörs direkt rätten till lika tillgång till utbildning .
Varför tiger kommissionen om detta ?
Vill den privatisera även utbildningen ?
Ekonomiska intressen ges mycket stort utrymme i avtalen , medan däremot offentliga intressen är mycket begränsade .
Det målas upp en bild av den fattige poeten .
Men här handlar det om ett fullständigt saluförande av Titanic soundtracks .
Dessutom har förhållandet mellan WIPO och TRIPS inte klarlagts , i synnerhet som delar av båda fördragen överlappar varandra .
Nu skulle man kunna säga : Ja det är klart , TRIPS , skillnaden är trade related intellectual property , men för WIPO handlar det ju huvudsakligen om handelsrelaterade aspekter .
Därför : Var är avgränsningen mellan de båda fördragen , och skall det finnas något samarbete ?
Om ja , i vilken form ?
Skall det med WIPO skapas ett precedensfall för att också fullständigt göra TRIPS underordnat EU : s ansvarsområde ?
Allt som allt finns det i förslaget fortfarande ett avsevärt behov av förklaring och förbättring .
Jag förväntar mig av kommissionen information om de frågor som ställts , för att jag överhuvud taget skall avge någon röstförklaring för min grupp .
Herr talman !
Ett tack till vår föredragande för det utmärkta betänkandet där hon likväl drar slutsatsen att vår anslutning till de båda WIPO-avtalen , i vår egenskap av gemenskap , inte bör inskränka sig till en liten institutionell förändring , hur viktig den än är , utan ge möjlighet åt Europeiska gemenskapen och WIPO-församlingen att arbeta tillsammans .
Ratificeringen är också nödvändig med tanke på utvidgningen av Europa .
Men bakom gemenskapens anslutning skönjs ett mål , som ännu är för virtuellt i mina ögon och ändå för offensivt i vissa medlemsstaters ögon .
Det handlar om att bekräfta en europeisk kulturpolitik om vilken jag väntar mig av oss , parlamentet , kommissionen och rådet , att vi är överens .
Om man säger kulturpolitik måste man säga försvar av skapandets roll , erkännande av upphovsmännen och framställning av en krävande kultur .
Och än mer nu då Europa skall införa en ny politik för upphovsrätt och närstående rättigheter är det brådskande - det har just betonats flera gånger - att fastställa och åter fastställa vad en upphovsman är .
Vi är i det avseendet ännu alltför vaga och de nya teknikerna kräver hädanefter att vi anstränger oss för att förtydliga detta .
Herr talman , ärade kommissionär !
Upprättandet av WIPO-avtalen utgjorde ett betydande positivt steg i utvecklingen mot ett globalt informationssamhälle .
Avtalen sammanfattar ett upphovsrättsligt arv från flera decennier och utgör en grundligt övervägd , välbalanserad lösning på frågan om reglering av upphovsrätt och närstående rättigheter .
Avtalens ikraftträdande och deras slutliga form beror utöver denna rekommendation dock även på parternas eget genomförande av dem .
I USA har WIPO-avtalet redan trätt i kraft med hjälp av Digital Millennium Corporate Act , och med detta lagstiftningsförfarande har man lyckats bevara den finkänsliga balansen i WIPO .
Också EU måste enligt överenskommelsen avancera i lagstiftningsarbetet inom WIPO .
Det är också oroväckande att det förra parlamentets ståndpunkter inte stödjer WIPO : s välbalanserade system .
Yttrandet om direktivet om upphovsrätt i den första behandlingen slog särskilt fel , och balansen är på väg att utvecklas i en ur europeisk synvinkel skadlig riktning .
De föreslagna rekommendationerna bidrar inte till att förbättra kulturens ställning i Europa , tvärtom .
De ändringar som parlamentet föreslagit skulle snarast göra det lättare för de etablerade mediaföretagen på marknaden att flytta över sina gamla , över 80-procentiga marknadsandelar till en ny miljö med osmidig och överdimensionerad upphovsrättsreglering .
Nu talar jag alltså inte om Charlotte Cederschiölds rekommendation , som är ett alldeles utmärkt dokument , utan om de upphovsrättsliga frågor som det förra parlamentet har behandlat .
Jag vill alldeles särskilt tacka fru Cederschiöld för att hon i sitt inlägg t.ex. har klargjort begreppet tillfällig kopia .
I WIPO-avtalet har man inte medvetet tagit ställning till tillfälliga kopior .
Om dessa tekniska kopior omfattades av skydd , skulle dataöverföringen - vilket alldeles riktigt konstateras i rekommendationen - bli dyr och komplicerad , utan någon anledning .
Det är ju fråga om samma situation som om brevbäraren var tvungen att betala upphovsrättsavgift då han leverar en bok till kunden som denne sedan läser .
Den verkliga fördelen med kultur är att konst och information säkert och enkelt kan föras över direkt från konstnären till användaren , konsumenten .
Den nya verksamhetsmiljön erbjuder först och främst ofantliga möjligheter att skapa och sprida kultur på ett helt annat sätt än någonsin tidigare .
Det är viktigt att alla parters intressen beaktas .
Detta har parlamentet velat beakta i sin egen rekommendation .
Herr talman !
På området skydd av upphovsrätten tycks verkligheten alltid ligga långt före bestämmelserna .
Utvecklingen av ekonomin , uppkomsten av nya kontraktsformer , de tekniska innovationerna är alla fenomen som innebär regelbundna och snabba förändringar som de ansvariga bör beakta vid utformandet av bestämmelserna .
På det området är processen för bestämmelsernas utformande en mekanism som rör sig långsamt , alldeles för långsamt i förhållande till de snabba förändringarna av den verklighet som de avser att reglera .
Om det påståendet stämmer i samtliga fall , är det ännu mer uppenbart när multinationella , överstatliga organ , som WIPO ( Världsorganisationen för den intellektuella äganderätten ) är involverade , där man har diskuterat de avtal som man avser att ändra .
När vi skall godkänna ratificeringen av dessa avtal , bör vi fråga oss om de motsvarar de mest aktuella behoven på området i fråga .
Svaret kommer knappast att bli positivt .
Det råder inga tvivel om att dessa avtal aktualiserar bestämmelserna på området , men det råder inte heller några tvivel om att det för närvarande är många problem som inte får någon lösning .
Encyclopedia Britannica har nyligen lagts ut på Internet och uppkomsten av virtuella bibliotek har uppenbarat att många problem återstår att lösa .
Den lösning som har valts av exempelvis ett av de främsta virtuella biblioteken - som tillhör mitt universitet , universitetet i Alicante - innebär att man utesluter verk med gällande upphovsrätt , och det hämmar i stor utsträckning utvecklingen av den här typen av virtuella bibliotek .
Å andra sidan kommer ratificeringen av avtalen att vara av ringa betydelse .
De problem som dessa löser har redan fått en god lösning i direktivet om harmonisering av vissa aspekter av upphovsrätt och närstående rättigheter i informationssamhället .
De flesta stater har redan antagit den lagstiftning som ligger till grund för de avtal som nu ratificeras .
Slutligen vill jag påpeka att de lagändringar som har införts i vissa länder , i Spanien till exempel , har inneburit en lösning på vissa konflikter , samtidigt som de har gett upphov till andra som är vanliga när det handlar om att prissätta rättigheter och material .
När man behandlar en så känslig fråga som denna bör man erbjuda lösningar som i lika utsträckning tar hänsyn till de intressen som står på spel .
Det är en förutsättning för att bestämmelserna skall kunna accepteras . .
( NL ) Herr talman !
Jag skulle gärna vilja börja med att gratulera föredraganden till det arbete hon lagt ner .
Kommissionen har intrycket av att hon arbetat snabbt och noggrant .
Det är viktigt .
Det passar sig för kommissionen att uttrycka sin tacksamhet till föredraganden .
För att direkt tala om kommissionens slutsatser : de överensstämmer med slutsatserna i förslaget till rekommendation .
Det betyder alltså att kommissionen instämmer i parlamentets ratificering .
Jag skulle gärna vilja betona båda avtalens betydelse .
WIPO-avtalet om upphovsrätt och WIPO-avtalet om utövande konstnärer och ljudupptagningar är båda två framsteg för ett internationellt immaterialrättsligt skydd och skydd av närstående rättigheter , och därmed är de en väsentlig förbättring av Bern- och Romkonventionerna .
De båda avtalen bidrar till en hög skyddsnivå för verk och andra saker , men de ger publiken tillgång till innehållet via elektroniska nät .
De två avtalen tillåter explicit att gemenskapen blir en fördragsslutande part och får en viktig uppgift när det gäller förvaltning på det här området .
Gemenskapens godkännande av avtalen har därför stor betydelse eftersom det visar att gemenskapen fäster stor vikt vid immaterialrätten .
Ett godkännande leder också till ett större internationellt erkännande av Europeiska unionens roll med avseende på upphovsrätt .
På internationell nivå finns det ett stort stöd för att avtalen skall träda i kraft snabbare .
De har nu ratificerats av tretton , respektive tolv , medlemsstater i WIPO , bland annat Förenta staterna .
Om de skall träda i kraft så snabbt beror till stor del på Europeiska unionen eftersom det behövs trettio ratificeringshandlingar för att avtalen skall träda i kraft och de handlingar som undertecknas av Europeiska unionen och medlemsstaterna samt av de associerade länderna är mycket viktiga för att komma upp i det antalet .
Även många utvecklingsländer förväntar sig att Europeiska unionen snabbt skall ratificera avtalen , det skulle nämligen vara en stark signal över hela världen .
Inom den ramen har parlamentet redan haft en mycket viktig roll vid diskussionerna om förslaget till direktiv om upphovsrätt i informationssamhället , vilka ledde till att Barzantibetänkandet godkändes i februari 1999 .
Det här direktivet är ett nödvändigt motstycke till det föreslagna beslutet och omfattar huvudsakligen de viktigaste principerna i WIPO-avtalen .
Europaparlamentet måste nu ännu en gång följa det särskilda samtyckesförfarandet enligt artikel 300.3 .
Den rätta signalen till yttervärlden , i form av den här rekommendationen , är av stor betydelse .
Kort sagt , för att åter upprepa kommissionens slutsatser : den stöder förslaget till rekommendation och hoppas att det skall ha stor betydelse för hela den värld som är intresserad av immaterialrätt .
Tack , herr kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
11.30 .
( Sammanträdet avslutades kl .
23.55 . )
