 
Parentation I går avled Bettino Craxi , före detta ledamot av Europaparlamentet , i Hammamet i Tunisien .
Bettino Craxi var ledamot av det här parlamentet från den 17 juli 1979 till den 20 augusti 1983 och från den 25 juli 1989 till den 30 april 1992 .
Craxi var också ordförande för rådet i sin egenskap av premiärminister för Republiken Italien , en post som han innehade från den 4 augusti 1984 och fram till sin avgång den 3 mars 1987 .
Får jag be er att hålla en tyst minut till hans minne .
( Parlamentet höll en tyst minut . )
 
Justering av protokollet från föregående sammanträde Protokollet från gårdagens sammanträdet har delats ut .
Finns det några synpunkter ?
Herr talman !
Jag skulle vilja ta upp en sak innan vi inleder fiskeridebatten .
De ärade ledamöterna känner kanske till den förfärliga tragedin med förlusten av en fiskebåt och hela besättningen på sju man i Skottland .
Solway Harvester sjönk med man och allt nära Isle of Man , när man fiskade efter musslor tidigare i år .
Besättningen på sju man kom från det lilla fiskesamhället Whithorn och kringliggande orter i Galloway i sydvästra Skottland .
Jag vet att jag talar för alla åtta parlamentsledamöterna från Skottland och för alla kolleger i denna kammare , när jag ber er att på Europaparlamentets vägnar sända ett kondoleansbrev till det skotska parlamentets talman , Donald Dewar .
Denna tragedi är kanske en läglig och ledsam påminnelse för oss alla , när vi påbörjar ytterligare en debatt om fiskeindustrin , om att tappra män och kvinnor varje dag riskerar sina liv i ett av de farligaste yrkena i världen för att skaffa fisk till våra bord .
Jag förlitar mig på att talmannen kommer att stödja denna begäran .
( Applåder ) Herr Stevenson !
Jag skall be ordföranden att skicka den här skrivelsen .
Det tycker jag verkar klart .
Herr talman !
I egenskap av ordförande i fiskeriutskottet och å mina kollegors vägnar vill jag solidarisera mig med vår kollega från Skottland , Stevenson , och den begäran han nyss lade fram .
Tyvärr har också vi nyligen haft ett olyckstillbud med en galicisk fiskebåt med galicisk och portugisisk besättning , Ros Alcedo , som började brinna i Gran Sol vatten .
Tyvärr är olyckshändelser av det här slaget betydligt vanligare än vad vi skulle önska , och därför vill jag påminna om att vårt utskott har begärt att få utarbeta ett initiativ till betänkande om orsaker bakom haverier och den fara yrkesfiskare löper .
Jag hoppas att betänkandet godkänns eftersom dessa hårt utsatta yrkesmän verkligen är i behov av kammarens och allas vårt stöd .
Tack , herr Varela .
 
Resultatet av de fleråriga utvecklingsprogrammen för fiskeflottorna ( 1997 ) Nästa punkt på föredragningslistan är betänkande ( A5-0096 / 1999 ) av Cunha för fiskeriutskottet om kommissionens årsrapport till rådet och Europaparlamentet om resultatet av de fleråriga utvecklingsprogrammen för fiskeflottorna vid utgången av 1997 ( KOM ( 1999 ) 175 - C5-0109 / 1999 - 1999 / 2112 ( COS ) ) .
Hudghton har begärt ordet i den här frågan .
Jag hoppas att ledamöterna uppskattar mitt starka intresse i denna fråga .
Jag vill , i enlighet med artikel 144 , väcka förslag om att Cunhas betänkande återförvisas till utskottet , och jag gör det med Verts / ALE-gruppens stöd .
I måndags framförde min kollega MacCormick tvivel om tillåtligheten för en del av punkt 6 i Cunhas betänkande , vilken inbegriper mycket känsliga frågor , som mycket väl kan komma upp igen i dag .
Men innan vi kommer dit , jag anser också att punkt 6 och förslagen däri omges av viktiga politiska och praktiska tvistefrågor .
Det skulle ligga i allas vårt intresse att försöka nå samstämmighet om vårt handlingssätt i denna fråga .
Därför skulle ytterligare diskussion i fiskeriutskottet , liksom även möjligheten att få ett yttrande från utskottet för rättsliga frågor och den inre marknaden , vara till stor hjälp för alla sidor i diskussionen .
Med tanke på de tvivel och vissa av de meningsskiljaktigheter som omger punkt 6 , skulle en återförvisning även möjliggöra och erbjuda ett tillfälle till ytterligare samråd , både med industrin och med våra sakkunniga i kommissionen och på annat håll .
Jag begär att vi röstar om att återförvisa betänkandet till utskottet och att vi åter tar upp det här i kammaren i sinom tid , efter ytterligare behandling .
Jag ber också om att denna omröstningar , om den genomförs , skall genomföras med namnupprop .
Herr Hudghton !
Ni gör mycket riktigt en formell begäran om återförvisning till fiskeriutskottet på grundval av artikel 144 i arbetsordningen .
Vi känner alla till de regler som gäller för detta .
Vid en sådan begäran kan en förespråkare och en motståndare ha ordet och även föredraganden eller utskottets ordförande om det behövs .
Finns det en förespråkare för denna nyss framlagda begäran ?
Herr talman !
Som Hudghton sade och som ledamöterna i kammaren nog kommer ihåg , bad jag i måndags om ordet för att säga att jag anser att en del i detta betänkande är otillåtligt , eftersom det saknar en rättslig grund .
Detta är snarast ett " domedags " vapen , och det skulle göra mig olycklig om vi tvingades använda det , när vi har en enklare metod att tillgå för att behandla ärendet på nytt , innan det slutligen kommer tillbaka till kammaren .
Det är en sak av högsta vikt .
I punkt 6 i Cunhas betänkande , som jag förstår den - och som många av mina kolleger förstår den - föreslås i själva verket en underminering av principen om relativ stabilitet som sedan 1983 har utgjort själva grunden för den gemensamma fiskeripolitiken , och som kommissionär Fischler under utfrågningen inför denna kammare faktiskt sade var av grundläggande betydelse för den gemensamma fiskeripolitiken .
Införandet av ett system för kvotbestraffningar skulle underminera den gemensamma politiken svårt , men det är just vad som föreslås i punkt 6 .
Betänkandet bör återförvisas till utskotten för behandling , både till fiskeriutskottet och till utskottet för rättsliga frågor och den inre marknaden .
Jag har nöjet att be kammaren att stödja Hudghtons förslag .
Herr talman !
Jag är emot det förslag som lagts fram .
Först och främst för att Cunhabetänkandet är ett betänkande som har godkänts av en majoritet i fiskeriutskottet .
Och inte bara det .
Den grundtanke som genomsyrar betänkandet är den som traditionellt sett parlamentet har fört fram i sina successiva betänkanden om utvärderingen av FUP ( flerårigt utvecklingsprogram inom fiskerisektorn ) .
För att besvara MacCormicks fråga om man i punkt 6 motsätter sig eller inte principen om relativ stabilitet , så vill jag säga att man i punkt 6 under inga omständigheter bestrider principen om relativ stabilitet .
Där föreslås bara , som en möjlig sanktion för dem som inte följer FUP , att de som mest förstör resurserna tillfälligt skall få sina kvoter indragna , det rör sig varken om en definitiv indragning eller om en överföring av kvoter från en medlemsstat till en annan .
Sammanfattningsvis kan man säga att principen om relativ stabilitet bevaras samtidigt som också sättet att använda sig av principen om relativ stabilitet bevaras , vilket många är rädda för .
Jag vidhåller därför att det inte finns någon som helst möjlighet att denna princip , denna heliga princip inom gemenskapsfisket , skall angripas .
Det är helt enkelt allvarliga sanktioner som föreslås - och eftersom de är kännbara klagar en del - för att effektivt värna om resurserna .
( Applåder ) Mycket kort skulle jag vilja säga att det inte handlar om principen om relativ stabilitet av det enkla skälet att det inte finns någon överföring av kvoter mellan medlemsstater , det handlar inte om det .
Vi talar dessutom om en tillfälligt avskaffande av kvoter för att tvinga medlemsstaterna att uppfylla målen i de fleråriga utvecklingsprogrammen .
Detta blir ännu klarare med ett godkännande av ändringsförslag 3 av Ford .
Jag vill , som föredragande , yrka på ett godkännande av detta .
För det andra vill jag säga att målet för punkt 6 i mitt betänkande är till för att just se till att Europeiska unionen skapar ett effektivt sanktionssystem , för om vi inte lyckas skapa sanktioner som tvingar länderna att uppfylla målen i de fleråriga utvecklingsprogrammen kommer de att bli meningslösa och vad värre är , bli ett instrument för diskriminering mellan de medlemsstater som uppfyller dem och minskar sina flottor och de som inte uppfyller dem och slipper sanktioner .
( Applåder ) Vi skall nu genomföra omröstningen om begäran om återförvisning till fiskeriutskottet .
Det är en omröstning med namnupprop .
( Begäran avslogs . )
Punkten kommer att stå kvar på föredragningslistan .
MacCormick har ordet .
Herr talman !
Artikel 143.1 : " När en debatt om en bestämd punkt på föredragningslistan inleds kan förslag väckas om att avvisa denna punkt som otillåtlig .
Ett sådant förslag skall omedelbart gå till omröstning . "
Jag väcker förslag om att avvisa punkten som otillåtlig och begär att ni omedelbart låter det gå till omröstning .
Jag blev verkligen inte imponerad av de argument som jag hörde tidigare .
Herr MacCormick !
Även här gäller regeln att en förespråkare och en motståndare kan få ordet .
Vem är för det här förslaget om att i enlighet med artikel 143 i arbetsordningen inte behandla denna punkt på föredragningslistan på grund av otillåtlighet .
Herr talman !
Jag kan gladeligen stödja min kollegas förslag om otillåtlighet , det vill säga otillåtligheten för punkt 6 i betänkandet .
Det finns tillräckliga tvivel om lagenligheten för förslaget som gäller automatiska kvotminskningar för en förklaring att punkt 6 - inte resten av betänkandet - är otillåtligt . )
Herr talman !
Det förvånar mig att en del ledamöter använder sig av samma argument som vid tidigare tillfällen , under föregående punkt togs nämligen också tillåtligheten för punkt 6 upp .
Jag tror att de flesta av oss ledamöter har klargjort att vi är för nämnda punkt och att vi redan har röstat om detta .
Vill ni så upprepar jag samma argument .
Punkt 6 strider inte mot principen om relativ stabilitet , principen respekteras och fördelningssättet respekteras .
Föregående talare säger sig vara tveksam .
Man måste känna sig säker för att kunna säga att man förkastar punkt 6 .
Är man tveksam måste man få det hela klargjort först .
Jag är inte tveksam , herr talman , och kammaren har redan visat detta .
Herr talman !
Med anledning av vad som här har sagts vill jag ta upp en annan ordningsfråga vad gäller arbetsordningens efterlevnad .
Vi har redan röstat om grunden .
Vi har redan röstat om huruvida en av de principer som tas upp i punkt 6 är tillåtlig eller inte .
En stor majoritet har förkastat ett återförvisande till utskott , vilket får mig att tolka detta som att punkten i fråga var tillåtlig .
Med detta ordklyveri kan vi inte än en gång rösta om samma fråga och säga att man nu skall tillämpa artikel 143 , eftersom man då anför samma skäl av otillåtlighet .
Jag menar att otillåtlighet tas upp i artikel 143 , otillåtlighet på grund av formella skäl .
Det stod inte med på föredragningslistan , det saknades vissa språkversioner etc . , men inte på grund av en fråga om grunden och än mindre om denna redan har diskuterats och lagts fram till omröstning .
Vi kan inte komma med ännu en ordningsfråga genom att använda oss av en annan artikel när kammaren redan har uttalat sig om grunden och sagt att man inte ämnar återlämna den till utskottet .
Nu får det vara nog med parlamentariskt ordklyveri .
Frågan bör avgöras precis som den redan har avgjorts av de flesta av oss som uttalat sig här i kammaren .
( Applåder ) Jag skall rekapitulera det hela .
Ett andra förslag har nu lagts fram i enlighet med en annan artikel i arbetsordningen och det måste jag som talman uppmärksamma .
Spelreglerna är klara .
En talare för och en talare mot har haft ordet och det har även utskottets ordförande .
Jag ger först ordet till föredraganden , Cunha , innan vi genomför omröstning med namnupprop .
Herr talman !
Jag skall inte tala för eller emot , jag vill bara säga att vi här är beskådar en fars .
Herr talman , var vänlig och läs arbetsordningen noga , för det vår kollega begärde har vi redan röstat om .
Det vore väldigt allvarligt om vi röstade enligt artikel 143 igen .
Detta är en oacceptabel fars !
( Applåder ) Herr talman !
Parlamentet har klart och tydligt uttalat sig i den här frågan och vi kan inte rösta två gånger om samma sak .
Jag vill uppmärksamma er på detta , det är nämligen en princip som vi alltid har respekterat .
Ordförandeskapets uppförande är just nu fullständigt oacceptabelt .
( Applåder ) Tyvärr , herr Barón Crespo !
Jag kan tänka mig hur ni känner er .
Det är emellertid inte helt rätt .
Nyss genomfördes en omröstning i enlighet med artikel 144 , det är återförvisningen till utskottet .
Den omröstningen har vi haft och återförvisningen förkastades .
Punkten står alltså kvar på föredragningslistan .
Vidare , och det kan ni inte klandra mig för , har ett andra förslag lagts fram , nämligen om att förklara ärendet otillåtligt .
Det är en annan artikel , artikel 143 i arbetsordningen .
( Förslaget förkastades . )
Herr talman och kära kolleger !
Europeiska kommissionens rapport om det första verksamhetsåret för det fjärde fleråriga utvecklingsprogrammet för fisket , det så kallade FUP IV för perioden 1997-2001 , visar att det 1997 skedde en minskning på 2 procent av gemenskapens flottkapacitet i bruttotonnage och 3 procent i maskinstyrka .
Härigenom var gemenskapsflottan den 1 januari 1998 nära 16 procent mindre än slutmålet för FUP IV när det gäller maskinstyrka och 7 procent när det gäller bruttotonnage .
Det finns några djupa förbehåll mot denna uppenbart optimistiska helhetsbedömning , av effektiviteten i de fleråriga utvecklingsprogrammen som instrument för att anpassa gemenskapsflottans storlek till tillgängliga fiskbestånd .
Det första förbehållet gäller svårigheterna att jämföra mål och avsikter mellan FUP III och FUP IV , på grund av att mätkriterierna och segmentindelningen av olika flottyper ändrats .
Det andra förbehållet vi har är att vi fortfarande har olika mätkriterier i varje medlemsstat , vilket gör utvärderingarna svåra att jämföra .
Jag måste för övrigt säga att kommissionen i sin rapport utfärdar en varning för just den bristande tillförlitligheten i de uppgifter som läggs fram .
Det tredje förbehållet vi har mot rapportens uppenbart optimistiska bedömning gäller det faktum att uppfyllandet av dessa mål är mycket olika mellan medlemsstaterna , där två inte uppfyller målen och en har lämnat information på ett oacceptabelt sätt .
I motsats till detta finns det medlemsstater , som exempelvis Portugal , Spanien , Danmark , Irland och Förenade kungariket , som redan har uppfyllt eller mer än väl uppfyllt de slutmål som fastställts i FUP IV - Portugal har mer än väl uppfyllt dem .
Till följd av detta föreslår jag främst två typer av åtgärder i mitt betänkande .
Den första typen av åtgärder består av att harmonisera mätkriterierna och segmentindelningen av flottorna och göra dem enhetliga , så att man kan göra komparativa , precisa och kontinuerliga bedömningar av gemenskapsflottan i varje medlemsstat .
Detta är grundläggande för att de fleråriga utvecklingsprogrammen skall vara effektiva .
Den andra typen av åtgärder handlar om behovet av gemensamma bestämmelser som framför allt innehåller ett effektivt sanktionssystem .
Därför , och bara därför , föreslår jag i mitt betänkande som exempel - jag vill betona det - att kvoterna skall upphävas för de medlemsstater som inte uppfyller målen för att tvinga dem att uppfylla dem .
Därför ansåg jag det vara lämpligt att acceptera ändringsförslag 13 av ledamoten Ford , för att understryka att detta upphävande är temporärt .
Jag vill understryka att det inte handlar om någon överföring av kvoter mellan medlemsstater , det handlar inte om någon kränkning av principen om den relativa staten , det handlar bara om ett temporärt upphävande för att politiskt tvinga länderna att uppfylla de fleråriga utvecklingsprogrammen .
Detta är mycket viktigt , eftersom de ekonomiska sanktionerna inom fonden för fiskets utveckling varit helt verkningslösa .
Om inte detta sker har inte medlemsstaterna några motiv att uppfylla de uppställda målen .
Om dessutom några uppfyller dem och andra inte och de som inte uppfyller dem slipper straff , bidrar vi faktiskt till en allvarlig diskriminering i tillämpningen av den gemensamma fiskeripolitiken mellan medlemsstater och vissa fiskare kommer att drabbas hårdare än andra .
Jag vill slutligen säga att om dessa två typer av åtgärder som föreslagits i mitt betänkande inte genomförs , kommer de fleråriga utvecklingsprogrammen för fisket inte bara vara verkningslösa , totalt verkningslösa , utan värre än så , de kommer ett vara ett element för diskriminering och snedvridning av konkurrensen mellan medlemsstater , mellan fartygsägare och mellan fiskare .
I så fall skulle det vara bättre att avskaffa dem .
( Applåder ) Herr talman !
Vi står ännu en gång inför kommissionens rapport om resultatet av de fleråriga utvecklingsprogrammen för fiskeflottorna denna gång för år 1997 .
Än en gång förvånas vi över hur kommissionen har kunnat basera en rapport på sådana meningslösa uppgifter som en del av medlemsländerna lämnat , något som enligt vår mening än en gång gör dokumentet i stort sett helt oanvändbart .
I rapporten kan man se att det finns fyra olika förhållningssätt när det gäller skyldigheten att följa det fleråriga utvecklingsprogrammet inom fiskerisektorn ( FUP ) .
Några få skickar , förutom att följa de allmänna målen att rekonstruera flottan , harmoniserade uppgifter - så som gemenskapsnormerna kräver - kan man tillägga .
Andra , de flesta , fortsätter att skicka in uppgifter där bruttotonnage ( BT ) och bruttoregisterton ( BRT ) blandas ihop , vilket gör det mycket svårt att kontrollera hur minskningen av tonnage uppfylls .
I den tredje gruppen finns två länder som under inga omständigheter uppfyller FUP : s allmänna mål .
Slutligen finns ett land som unnar sig lyxen att inte skicka in en enda uppgift , något som man har gjort tre år i rad .
Detta är inte bara en oacceptabel diskriminering av de länder som uppfyller de allmänna målen genom att utsätta sina flottor för stora uppoffringar , utan också för dem som inte uppfyller målen , men som åtminstone fullgör sin skyldighet att lämna in uppgifter , skyldigheter som de straffbeläggs för att inte fullgöra .
För ett medlemsland , som genom att vända ryggen till gemenskapens regelverk tre år i rad har dolt sina uppgifter , kommer detta inte att inträffa , och eftersom man inte känner till dess siffror kan man inte heller straffbelägga landet i fråga .
Detta är ett så stort lurendrejeri att vi enbart med stor ansvarskänsla kan uppmuntra de länder som fullgör sina skyldigheter att fortsätta anpassa sina flottor till nuvarande resurser och inte tvärtom .
Det tråkiga är att vi fortsätter att ålägga skyldigheter när vi i dagens läge inte ens vet hur många båtar och hur stort tonnage som finns i gemenskapsflottan .
Med anledning av detta har kommissionen informerat om att det nästkommande månad kommer att finnas en expertstudie tillgänglig om hur stora medlemsländernas flottor är utom för ett land , och jag skulle vilja veta om det är samma land som alltid .
Innebär detta att Cunha för varje år måste lägga fram ett av sina utmärkta betänkanden om hur FUP uppfylls samtidigt som han på nytt måste varna för faran om några av medlemsländerna fortsätter att tro att bevarandet av gemenskapsresurserna alltid faller på någon annans bord ?
Herr talman , det måste bli ett stopp på detta .
Därför är vår föredragandes begäran om att sanktioner skall införas i form av minskade fiskekvoter , inte bara för dem som inte fullgör sina skyldigheter utan också för dem som envist framhärdar bakom ockultism och bedrägeri , en väl genomtänkt begäran .
De påföljder som finns medtagna i det nya finansiella instrumentet för utveckling av fisket ( FIUF ) är mycket riktigt ett steg i rätt riktning , men inte tillräckligt för att förhindra alltför långvarig uraktlåtenhet .
Därför stöder vi föredraganden och dennes begäran om reellt stävjande åtgärder och vi anser , tvärtemot vad vissa andra tycker , att den här typen av straff är synnerligen rimliga .
För det första för att man nått den punkt där man måste slå där det gör som ondast .
För det andra för att även om kvoterna inte inkluderas i den strukturella politiken så är en bristande fullgörelse av FUP ett hot mot detta medel .
Det slutliga målet med gemenskapens fiskeripolitik är ju att skydda bestånden .
Herr talman , efter det som inträffade i morse vill jag säga en sak : Även om jag alltid har varit övertygad om att Cunhas betänkanden och förslag i den här frågan varit bra , så är jag än mera övertygad nu , jag tror faktiskt att han har satt fingret på den ömma punkten .
Jag hoppas att de andra två institutionerna som måste fatta ett beslut i frågan förstod att en tillämpning av effektiva sanktioner skulle kunna lösa problemet med en alltför stor gemenskapsflotta , vilket vi nu har , och att vi därmed skulle kunna värna om våra resurser och framför allt om våra fiskare .
Herr talman , ärade kollegor !
Den gemensamma fiskeripolitiken ser jag i huvudsak som en samling regler som alla aktörer måste följa .
Föreställ er ett parti schack där en spelare flyttar löparna diagonalt - enligt reglerna - men använder hästarna som om de vore torn och som dessutom försöker fortsätta att spela trots att han försatts i " schackmatt " .
Föreställ er dessutom att domaren tittar åt ett annat håll .
Detta är enligt min mening vad den föregående kommissionen gjorde .
Vi förlitar oss nu på att den nuvarande fullföljer sitt uppdrag som fördragets väktare och inte tillåter att " så många mål görs " .
Bevarandet av våra fiskeresurser är mycket riktigt avhängigt respekten för de avtal som fastställts när det gäller total tillåten fångstmängd ( TAC ) , kvoter , viloperioder samt ländernas åtaganden för att minska sina respektive flottor .
Om någon från detta sköra kortslott som vi tillsammans har byggt tar bort ett enda kort så rasar , ärade kollegor , hela konstruktionen .
Att följa FUP är ett absolut krav för att säkra jämvikten mellan resurserna och flottans kapacitet .
De olika medlemsländernas grad av fullgörelse när det gäller förpliktelserna mot FUP är som skillnaden mellan natt och dag , vilket betänkandet klart och tydligt visar .
I detta första betänkande finner vi länder som med stor ekonomisk och social kraftansträngning och med stora påfrestningar för sina respektive fiskeflottor och folk på ett korrekt sätt har fullföljt sina åtaganden .
Detta erkänns av såväl kommissionen som av Cunha i dennes betänkande .
Cunha , som jag tackar för ett utmärkt betänkande , förklarar också hur en del medlemsländer brister i sin fullgörelse samtidigt som han anger en bristande vilja hos några andra som dessutom vägrar att tillhandahålla tillförlitliga uppgifter .
Som föredraganden säger , så är det ofattbart att kommissionen har tolererat att ett land under så många år har underlåtit att lämna tillförlitlig information om sin flotta .
Något som förmodligen var möjligt tack vare den dåvarande kommissionens politiska svaghet .
Det finns dock andra skäl som jag skulle vilja ta upp och som ankommer på Europeiska kommissionen och medlemsländerna , det är nämligen nödvändigt att båda i den här nya etappen anstränger sig för att harmonisera de referenskriterier som skall gälla för att mäta tonnage och fartygens kraft .
Bara på det här sättet kan vi undvika att några gäckar reglerna , vilket är vad som sker nu .
Kommissionen måste , som Cunha säger i sitt betänkande , vara mera strikt när det gäller kriterierna för en segmentering av de nationella flottorna , man måste på ett bättre sätt fastställa de geografiska zonerna samt använda sig av sin sanktionerande kapacitet , må vara temporärt , för att förmå länderna att fullgöra sina åtaganden när det gäller att minska sina flottor .
Vi socialdemokrater kräver att kommissionen här i parlamentet lovar att man inte längre kommer att tolerera att FUP inte följs och att vissa länders bristande öppenhet inte heller kommer att tolereras , ett uppförande som bara skadar andra som gör allt för att försöka nå de mål som uppställts av FUP .
Kommissionen skall vid utövandet av sin behörighet se till gemenskapens bästa .
Herr talman !
Låt mig inledningsvis gratulera Cunha till ett lysande betänkande som vi i det stora hela kan stödja .
Vi ser allvarligt på kommissionens anmärkningar i årsrapporten om resultaten av de fleråriga utvecklingsprogrammen för fiskeflottorna i gemenskapen .
Man bör också notera att rapporten är från 1997 och att vi i dag skriver 2000 .
Årsrapporten präglas av en rad ändringar i referensgrunden och därmed komplicerade utvärderingar rörande mätningarna , som blir ännu svagare eftersom inte alla medlemsstater följer programmen .
Vissa länder uppfyller de slutliga målsättningarna för FUP IV och andra länder är mer eller mindre försenade .
Man talar dessutom om att det inte finns tillförlitliga uppgifter från andra länder .
Det är viktigt att påpeka att det kanske finns stora brister , eftersom det inte existerar några enhetliga jämförelsekriterier .
Cunha hänvisar i sitt betänkande till att målet med de fleråriga utvecklingsprogrammen är att skapa balans mellan de tillgängliga fiskeresurserna och den gemensamma fiskeflottans insats .
Det betonas att en väsentlig minskning av fiskeflottan är en förutsättning för att säkerställa en hållbar utveckling inom sektorn .
Här tänker jag inte minst på de unga som skall starta verksamhet .
Jag tänker på investeringar i nya fartyg .
Det är också en given förutsättning att de socioekonomiska offren skall fördelas på ett rättvist sätt mellan medlemsstaterna .
Vi är bekymrade över att en mängd medlemsstater är försumliga - ja , nästan likgiltiga - när de gäller att inrapportera pålitliga uppgifter om sin fiskeflottas status .
Det är dessutom mycket tydligt att det från en rad medlemsstaters sida bara visas ett litet intresse av att minska fiskeflottans kapacitet i enlighet med programmens målsättningar och beslut .
Fiskeriutskottet uppmanar kommissionen och medlemsstaterna att anta enhetliga och jämförelsebara kriterier för mätningar , och det måste vara ett absolut krav .
Kommissionen uppmanas vidare att öka kontrollen av utvecklingen inom medlemsstaternas flottor .
Detta stöder vi också fullständigt .
I förlängningen av den skärpta kontrollen uppmanas kommissionen att vidta och i givet fall skärpa åtgärder den redan vidtagit , för att tvinga medlemsstaterna till att uppfylla bestämmelserna om en reduktion av fiskeflottan .
Det kan ske i form av avslag till stöd för förnyelse och modernisering av fiskeflottan och i form av rättslig prövning vid EG-domstolen .
Cunha föreslår att medlemsstaternas bristande inrapportering av uppgifter kan medföra en minskning av fiskekvoterna .
Vi menar att detta inte är rätt väg att gå , eftersom vi inte anser att yrkesfiskarna skall straffas på grund av att medlemsstaterna är försumliga .
Vi har bett om delad omröstning om detta ändringsförslag .
Vi har också gjort detta i samband med hänvisningen till relativ stabilitet , eftersom vi menar att man här blandar ihop frågorna på ett sätt som kan riskera att snedvrida den princip som fastställs i fördraget .
För att sätta in den här debatten i sitt sammanhang , låt oss komma ihåg att det nuvarande fleråriga utvecklingsprogrammet för fiske ( MAGP ) , den fjärde generationen , inte alls följer de vetenskapliga råden från Lassenkommittén .
Kommittén rekommenderade stora minskningar av EU : s flottor , för att ge bestånden en chans att återhämta sig .
Rådet kunde inte godta det , så i den slutgiltiga förordningen föreskrivs relativt blygsamma minskningar .
Man avser minska EU : s totala flotta med endast 2,3 procent vad beträffar tonnage och 3 procent vad beträffar motorkraft under de fem år som programmet varar .
Som framgår av kommissionens rapport , var EU : s sammanlagda flottor i början av 1998 , bara ett år in i programmet , redan lågt under dessa mål .
Snarare än att visa hur duktiga medlemsstaterna har varit , visar detta i själva verket att de begärda minskningarna verkligen var mycket blygsamma och långt mindre än vad som var nödvändigt .
Icke desto mindre , och detta är den verkliga tvistepunkten , har många medlemsstater inte följt förordningen , och många av flottorna är för stora .
Vad gör man med dessa medlemsstater som sätter sig själva över gemenskapslagstiftningen och ignorerar sina åtaganden ?
Kommissionen har föreslagit flera saker : Den kan hålla inne strukturfonder , men det är ett effektivt verktyg bara om medlemsstaten verkligen använder fonderna .
Den kan dra medlemsstaten inför domstol , men det är tidsödande , dyrt och besvärligt .
I sitt förslag om den nyligen genomförda förnyelsen av FIUF föreslog kommissionen att medlemsstater som inte rättade sig skulle nekas tillgång till fisketillstånd enligt fiskeavtal med tredje länder .
Som man kunde vänta sig , vägrade rådet .
Vi måste finna medel som är effektiva för att övertala eller tvinga medlemsstater att respektera sina juridiska åtaganden .
Cunha bad kommissionen att överväga möjligheten till kvotsanktioner , om MAGP-målen inte respekteras .
Somliga anser att detta är ett brott mot principen om relativ stabilitet , men låt oss komma ihåg att principen om relativ stabilitet bara är en av principerna i den gemensamma fiskeripolitiken .
I den grundläggande förordningen sägs också att gemenskapens förvaltningssystem måste göra det möjligt att skapa en balans på permanent basis mellan resurser och utnyttjande .
Med andra ord , om alla bestånd havererar , är relativ stabilitet av en nollkvot inte värt särskilt mycket .
Vi tycker att idén åtminstone förtjänar ett seriöst övervägande .
Det finns redan ett tidigare fall i förordning 847 / 96 om de fleråriga tillåtna totalfångsterna .
Principen i förordningen är den , att om en medlemsstat överskrider sin kvot för vissa arter , minskas dess kvot för följande år , inte bara med den överfiskade mängden , utan med en extra mängd , som ökar ju större överfiskning har varit .
Detta är helt klart ett straff , men det ansågs inte vara ett brott av den relativa stabiliteten .
Cunhas uppslag kunde kanske ha varit mer omsorgsfullt formulerat , för att klargöra att ingen minskning skulle vara permanent , utan av begränsad varaktighet , och det är av den anledningen som vi kommer att stödja ändringsförslaget från PSE på denna punkt om att inkludera " temporärt " .
Jag är övertygad om att alla håller med mig om att vi måste finna sätt att se till att medlemsstaterna följer lagstiftningen .
Herr talman !
Analysen av det första tillämpningsåret för den fjärde generationens fleråriga utvecklingsprogram , som kommissionen har genomfört , visar att situationen ser mycket olika ut i de olika medlemsstaterna .
Medan några länder inte uppfyller de fastslagna målen eller inte lägger fram tillförlitliga uppgifter , finns det andra länder som inte bar uppfyller dem utan till och med går längre än de angivna målen , vilket är fallet med Portugal .
Gemenskapsflottan var således i början av 1998 mindre än slutmålet för FUP IV när det gäller maskinstyrka ( 16 procent mindre ) , och när det gäller bruttotonnage ( 7 procent mindre ) .
Men när det gäller Frankrike och Nederländerna har de ännu inte uppnått målen i FUP och för Italien känner man inte till några uppgifter .
Portugal har inte bara gått längre än det europeiska genomsnittet , med en minskning av 38 procent för tonnaget och 21 procent för maskinstyrkan , utan är det land som har minska sin flottas fiskeansträngningar mest , med allt vad detta innebär i förstörelse av fartyg , förlust av arbetstillfällen och hot mot nära 180 viktiga samhällens överlevnad .
Det finns alltså en klar obalans i Europeiska unionens fiskesituation , även om vi tillämpar den försiktighet som är nödvändig vid analys av de uppgifter som har lagts fram i rapporten , vilket föredraganden påpekar .
För Portugal är den aktuella situationen särskilt allvarlig och är i grunden ett resultat av en gemensam fiskeripolitik som inte tar hänsyn till särdragen i varje medlemsstat , även om det också ligger ett ansvar i den nationella politiken hos den som vill vara bästa eleven i uppfyllandet av de europeiska bestämmelserna .
Det står i dag klart att en fiskeripolitik som grundas på ett litet stöd till modernisering och förnyelse av flottan , på åtgärder för att förstöra fartyg och upphöra med verksamheten , på dåliga arbetsvillkor och låga löner för fiskarna , tillsammans med en stark yttre konkurrens , har bidragit till att drastiskt minska landets fiskekapacitet och håller på att framkalla en emigration av de portugisiska fiskarna till flottor i andra länder , främst till dem som inte har uppfyllt målen i de fleråriga utvecklingsprogrammen utan till och med har ökat sin fiskekapacitet .
Det är alltså nödvändigt med en långtgående förändring av den gemensamma fiskeripolitiken , och inte bara i den konkreta frågan om de fleråriga utvecklingsprogrammen , med speciell uppmärksamhet på särarten hos varje land , med speciella stöd till förnyelse och modernisering av flottan i medlemsstater som redan har uppfyllt målen , med stödåtgärder för att fiskesamhällena skall överleva , med en förbättring av fiskarnas livs- och arbetsvillkor och fastställandet av kompensationsbidrag vid förbudsperioder , vilket är fallet med sardiner i Portugal , eller vid eventuella andra nödvändiga minskningar av fiskeperioden .
Herr talman !
Införandet av det fjärde fleråriga utvecklingsprogrammet inom fiskerisektorn är synnerligen svårt .
Denna sektor har ju redan gjort avsevärda ansträngningar för att anpassa sin flottas kapacitet under de tidigare planerna .
Och ändå begär kommissionen att de skall fortsätta med kapacitetsminskningen .
Bortom en viss tröskel är emellertid inte flottans nivå tillräcklig för att hamn- och handelsinfrastrukturerna skall amorteras och vara lönsamma , vilket riskerar att leda till fullständigt oberättigade omlokaliseringar och minskningar av antalet båtar om vi behåller fångstkvoterna .
De utvecklingsplaner som utformats såsom planer för fortsatt minskning av flottan får således inte bli permanenta komponenter i den gemensamma fiskeripolitiken .
Därför kan inte ledamöterna av Gruppen Unionen för nationernas Europa godkänna betänkandet Cunha i dess nuvarande skick .
Därför har vår kollega Dominique Souchet ingett fem ändringsförslag som syftar till att påminna om att fångstkapaciteten bör anpassas och inte tvunget , systematiskt och ständigt minskas .
Vårt mål är nämligen att säkra att EU : s medlemsstaters fiskeflotta överlever .
Våra ändringsförslag anger också att det är svårt att genomföra en jämförelse mellan den tredje och fjärde planen på grund av att nya faktorer tillkommit , såsom fångsternas sammansättning och motorernas natur .
De påminner också om att det är svårt för medlemsstaterna att med kort varsel lämna de detaljerade och mångtaliga uppgifter som begärs av dem .
Vår grupp kommer dessutom att vara emot punkt 6 i resolutionsförslaget .
Det är nämligen inte Europaparlamentets sak att begära att de tillämpliga straffavgifterna i händelse av att planerna eller anmälningsförfarandena inte följs skall kunna bestå av ytterligare kvotminskningar .
Enligt vår åsikt finns det först och främst ingen rättslig grund för det och utvecklingsplanernas natur får hur som helst inte förändras .
Jag upprepar att deras syfte inte är att fiskeriverksamheten i Europa skall försvinna utan tvärtom att den skall kontrolleras för att säkra dess överlevnad .
Mot bakgrund av oljeutsläppet i Frankrike nyligen har vår grupp också ingett två ändringsförslag enligt vilka begärs att tillämpningen av minskningsplanerna skall låsas i de drabbade områdena .
Europaparlamentet i sin helhet upprördes ju i veckan av denna katastrof .
I vår grupp befann sig Dominique Souchet och Philippe de Villiers i katastrofens centrum i Vendée och rapporterade till oss hur brådskande det var att vidta solidaritetsåtgärder .
Det är uppenbart att fiskeriverksamheten i de drabbade områdena försvagas under en viss period .
Att på under sådana omständigheter vilja tillämpa restriktiva åtgärder på ett enhetligt sätt i Europeiska unionen utan att ta hänsyn till exceptionella situationer skulle kunna leda till ytterligare katastrofer .
Herr talman !
Mitt partis policy är att motarbeta den gemensamma fiskeripolitiken , eftersom vi anser att fiskeresurserna bör förvaltas av de individuella medlemsstaterna ensamma .
Följaktligen är jag också emot det fleråriga utvecklingsprogrammet ( FUP / MAGP ) , eller " skatan " , som vi kallar det i UK , den välbekanta svarta och vita fågeln som är så duktig på att urskillningslöst döda ungfåglar och som även är en berömd tjuv - vilket i mångt och mycket i Förenade kungariket är fiskeindustrins bild av den gemensamma fiskeripolitiken .
Men även om jag inte var emot det av allmänna skäl , skulle jag vara emot Cunhas betänkande på grund av dess specifika innehåll .
Den främsta anledningen till att jag är det härrör från formuleringar i rapporten , som till exempel i punkt a på sidan 4 , där följande formulering återfinns : " En lämplig politik för att bevara resurser är ett nödvändigt krav för att garantera framtiden för en lönsam och konkurrenskraftig fiskerisektor i gemenskapen . "
Om man betonar ordet " lämplig " , är mitt problem att " skatan " inte är en lämplig politik för att bevara resurser .
Från ett brittiskt perspektiv är den centrala bristen att vi har varit tvungna att acceptera ett stort antal utländska trålare i våra vatten , över vilka vi inte har någon direkt kontroll .
För oss handlar inte frågan om att för många båtar jagar för få fiskar , som kommissionen vill få oss att tro , utan om att för många EU-båtar jagar för få fiskar .
En mer grundläggande brist är kvotsystemet .
De senaste uppskattningarna är att 3,7 miljoner ton fisk kastas tillbaka döda varje år .
Detta är en verklig miljökatastrof .
Vi måste angripa kvotsystemet .
Det har varit helt och hållet verkningslöst vad gäller att kontrollera fiskeresurserna på något som helst sätt .
Jag kommer att rösta emot detta betänkande av Cunha , eftersom det skapar ännu fler sanktioner .
Det gör ännu fler fiskare till brottslingar .
Herr talman , fru kommissionär , ärade kollegor !
Jag tycker verkligen att det betänkande som utarbetats av föredragande Cunha är ett utmärkt betänkande , ett betänkande som kommer mycket lägligt , vilket var uppenbart i morse .
Jag tackar honom uppriktigt för detta .
Jag skall fatta mig kort .
Vi talar hela tiden om det rådande problemet mellan fiskeflottans storlek och befintliga fiskeresurser .
Vi talar om överkapacitet när det gäller fiske , överexploatering av resurser på grund av en överdimensionerad flotta .
Kommissionen igångsatte de så kallade fleråriga utvecklingsprogrammen inom fiskerisektorn ( FUP ) för att försöka få till stånd en jämvikt i nämnda relation .
Något som har visat sig är att FUP respekteras olika i olika länder .
En del har följt programmet till punkt och pricka med en minskning av sin flotta med upp till 40 procent , andra har inte uppfyllt några krav alls .
En del vägrar till och med att lämna uppgifter om hur programmet följs , och det allvarligaste av allt är att de som brister i sin fullgörelse också gör anspråk på att bli behandlade på samma sätt som dem som hårdnackat och smärtsamt har minskat sin fiskekapacitet med en påföljande ekonomisk och social uppoffring .
Därför är Cunhas betänkande viktigt och opportunt .
Här visar man kommissionen vilka de grundläggande problemen är : Projekt som är föga rigorösa , ojämn kontroll och framför allt bristande enhetlighet i de olika ländernas kriterier för att mäta sin flottas storlek .
Som om detta inte vore tillräckligt så informeras man i betänkandet om att effektiva påföljder för dem som brister i sin fullgörelse inte finns , något som till syvende och sist innebär att de mekanismer som skulle kunna vara användbara för det ändamål de skapades inte tjänar något till .
Därför måste kriterierna harmoniseras och vi måste effektivt bestraffa dem som inte fullgör sina åtaganden .
I Cunhabetänkandet nämns som exempel en minskning eller indragning - åtminstone temporär , om Fordbetänkandet godkänns - av kvoterna för det land som begått överträdelsen i fråga .
Vi får hoppas att parlamentet under plenarsammanträdet godkänner betänkandet , precis som det godkänts i fiskeriutskottet med de ändringsförslag föredraganden har hänvisat till , och att kommissionen och rådet verkligen noterar detta så att de kan ge ny styrka åt nyckelinstrumentet för att nå målen i gemenskapens nuvarande fiskeripolitik , det vill säga mål som baseras på en hållbar utveckling inom sektorn , vilket är vad vi från fiskeriutskottet vill se .
Herr talman !
Jag vill göra en grundläggande kommentar om Cunhas betänkande .
Jag har en viss förståelse för de politiska synpunkter som våra nationalistiska kolleger framförde i morse avseende punkt 6 , men vad beträffar deras sätt att ta itu med denna punkt , valde de fel tillvägagångssätt .
Det är inte lämpligt , och i omröstningen kom vi fram till att inte återförvisa betänkandet till utskottet .
Vi stöder inte heller åsikten att punkt 6 är otillåtlig .
Det bästa tillvägagångssättet är att rösta om betänkandet och följa den politiska logiken .
Jag har lagt fram ett ändringsförslag i vilket " temporärt avlägsnande av kvoter " ersätter antydningen i punkt 6 om att det skulle vara " permanent " , om medlemsstaterna inte följer bestämmelserna .
Om detta ändringsförslag , eller något likvärdigt , går igenom , kommer vi att stödja betänkandet .
Om inte , kommer vi att rösta emot det .
Ett sådant ändringsförslag kommer att sätta press på regeringarna att följa lagen , utan att man ger avkall på principen om relativ stabilitet , vilken , som vi alla mycket väl vet , har utgjort grunden i den gemensamma fiskeripolitiken sedan 1983 .
Detta är det bästa tillvägagångssättet , som vi också kommer att följa , och vi hoppas att de andra politiska grupperna kommer att tillåta att betänkandet går igenom med de nödvändiga ändringarna .
Herr talman !
Jag har två invändningar mot punkt 6 i Cunhas betänkande , vilket jag gratulerar honom till som helhet .
För det första , angående den automatiska minskningen av kvoter för medlemsstater som bryter mot bestämmelserna .
Min invändning är att följden av detta faktiskt är att sanktionerna missar sitt mål .
Om vi minskar kvoterna , är det fiskare och deras levebröd som kommer att drabbas .
Det är helt tvärt emot rättvisans principer att straffa vissa människor för andras fel .
Min andra invändning gäller hänvisningen till principen om relativ stabilitet .
I mina ögon är argumentet att punkten faktiskt undergräver denna princip övertygande .
I dess nuvarande formulering finns det i punkten en hänvisning till en automatisk minskning av kvoter , utan någon specificering beträffande omfattning eller tidsgränser .
Detta skulle kunna leda till en kraftig urholkning av traditionella fiskerättigheter .
Det är någonting helt annat än minskningar vid överfiskning , som ju helt enkelt återställer balansen .
Jag känner till ändringsförslaget i vilket det föreslås att minskningarna endast bör vara temporära , men jag anser att det skulle vara långt säkrare att ta bort hänvisningarna till kvoter och till principen om relativ stabilitet helt och hållet .
Jag inser fullständigt att vi behöver seriösa och effektiva straff , men vi måste se till att de respekterar den gemensamma fiskeripolitikens principer och drabbar dem som förtjänar dem .
Herr talman !
Cunhas betänkande är betydelsefullt , eftersom Cunha i betänkandet försöker undersöka hur medlemsstaterna uppfyller sina förpliktelser .
Om man inom Europeiska unionen enas om regler och bestämmelser , har medlemsstaterna och regeringarna självklart ett ansvar att rätta sig efter dessa .
Jag har inte några som helst svårigheter att stödja den principen , men hur skall en försumlig part bestraffas ?
Finns det i det här fallet ett behov av nya sanktioner ?
Om svaret är ja , är det då troligt att de sanktioner som föreslås av Cunha är effektiva ?
I punkt 6 försöker man ta itu med frågan om kvotsanktioner , som Cunha och Fraga Estévez stöder så helhjärtat .
Jag ber inte om ursäkt för att jag tog upp ordningsfrågor om detta ärende tidigare i förmiddags .
Det är tveksamt om förslaget om att använda automatiska kvotnedskärningar är lagenligt , det är opraktiskt och snudd på ogenomförbart , och det straffar fiskarna - inte medlemsstaterna - , vilket min skotska kollega påpekade för en liten stund sedan ; och viktigast av allt är att det hotar att undergräva principen om relativ stabilitet .
Fraga Estévez har helt riktigt påmint oss om att kvotstraff har tagits upp i detta sammanhang i tidigare debatter här i kammaren .
1998 debatterades ett liknande förslag , och det kan till och med ha haft samma upphovsman .
Den dåvarande kommissionären , Bonino , sade i sitt svar på debatten , och jag citerar : " Ett ändringsförslag innehåller förslag om sanktioner .
Kommissionen kan av flera anledningar inte godta detta förslag .
För det första eftersom automatiska minskningar av kvoterna för länder som inte fogar sig allvarligt undergräver den grundläggande principen i den gemensamma fiskeripolitiken , som är principen om relativ stabilitet . "
Hon sammanfattade genom att säga - jag citerar igen : " Jag skulle därför vilja be parlamentet om att på nytt överväga kvotminskningar som en sanktion , med tanke på dessa möjliga konsekvenser . "
Jag hoppas att den nya kommissionen kommer att slå in på samma linje efter dagens debatt .
Det är synd att Fischler inte är här och kan tala för sig själv , även om han , vid utfrågningen , gjorde mycket positiva kommentarer om relativ stabilitet , vilket jag välkomnar .
Det har lagts fram ändringsförslag för punkt 6 , men jag kan inte stödja dem , eftersom man i båda godtar principen om att använda kvotminskningar som ett straff .
Fastställandet av kvoter bör uteslutande baseras på vetenskapliga mål och på bevarandemål , inte användas som ett automatiskt straff .
Om försumliga medlemsstater skall uppmuntras till att uppfylla FUP-målen , måste ett effektivt sanktionssystem riktas mot regeringarna - inte mot fiskarna .
Vi har begärt delade omröstningar om punkt 6 , och jag hoppas att vi kommer att få möjlighet att utöva dessa , och jag hoppas att ledamöterna i denna kammare i princip kommer att motsätta sig användningen av kvotstraff som avskräckningsvapen i detta ärende .
Herr talman !
I den här debatten om de fleråriga utvecklingsprogrammen måste vi ha helt klart för oss vad slutmålet egentligen är .
Egentligen handlar det ändå om att skydda fiskbeståndet genom att begränsa fångsterna .
För att göra det möjligt för den här sektorn att följa kvoterna så har Europeiska unionen som kompletterande åtgärd givit medlemsstaterna i uppdrag att minska sina flottor .
De fleråriga utvecklingsprogrammen är alltså inget självändamål utan instrument för kvotregleringen .
Tyvärr måste jag konstatera att föredraganden vänder på mål och medel .
Det märks när han yrkar för att införa en kvotminskning för en medlemsstat som inte uppfyller de fleråriga utvecklingsprogrammen , oavsett om den respekterar kvoten eller inte .
På det sättet utropar han de fleråriga utvecklingsprogrammen till det högsta målet och degraderar kvoterna till praktiska instrument .
Medlemsstater som inte helt efterlever de fleråriga utvecklingsprogrammen men som respekterar kvoterna - vilket väl ändå är själva slutmålet - straffas orättvist hårt på det sättet .
Jag tänker i det fallet på Nederländerna som visserligen inte minskat sin flotta i så stor omfattning men som ändå med hjälp av en reglering av antalet dagar till havs , lyckas klara sig inom kvoterna .
Vore det inte rättvisare att ålägga de medlemsstater som ständigt överskrider sina kvoter , och alltså verkligen utgör ett hot för fiskebestånden , en extra minskning av fiskeflottan ?
Avslutningsvis förekommer starka tvivel angående de olika medlemsstaternas flottkapacitet .
Politik som grundar sig på otillförlitliga uppgifter är en dålig politik och skadar myndigheternas auktoritet .
Därför uppmanar jag kommissionen att snarast grundligt kontrollera medlemsstaternas uppgifter genom en sakkunnig och oberoende organisation .
Herr talman !
Först av allt vill jag tacka Cunha för hans stora sakkunskap .
Jag måste konstatera att han på ett bra sätt har klargjort ett antal fakta angående de fleråriga utvecklingsprogrammen .
Han har med rätta sagt att många uppgifter inte är tillförlitliga , att det är svårt att få fram de rätta uppgifterna och att det är ett av problemen med den europeiska fiskeripolitiken .
Så långt hyser jag alltså stor uppskattning för det hela .
Min kritik gäller några andra punkter .
Om man nämligen konstaterar att uppgifter inte är tillförlitliga , att ett program egentligen är ett kompletterande program och vidare yrkar för sanktioner som är mycket långtgående , då kan det leda till diskriminering av medlemsstater och absolut av fiskare .
När man konstaterar att uppgifter inte är tillförlitliga så måste man också se till de sanktioner som hanteras .
Annars skulle det kunna hända att länder som inte helt uppfyller en del av utvecklingsprogrammen och som redan straffas ekonomiskt för det - det är ju faktiskt så i den politik som redan förs - sedan straffas en gång till medan länder som inte lämnar lika fullständiga uppgifter går fria .
Det får inte vara på det sättet , tycker jag .
Jag skulle också vilja yrka för , även det inom ramen för det här betänkandet , att vi hittar ett bättre sätt att jämföra uppgifter mot varandra i Europeiska unionen .
Harmonisering av uppgifter , bättre kontroll och en riktad politik på grundval av det .
En annan punkt som jag skulle vilja yrka för i det här sammanhanget är att de sanktioner som görs begränsas till den politik som förs .
I det här fallet till de fleråriga utvecklingsprogrammen och det innebär att medlemsstater som på ett eller annat sätt inte helt kan uppfylla dem eventuellt kan utsättas för sanktioner i just det avseendet .
Det betyder att de kan få mindre pengar .
Det är en sanktion som hör till den här politiken och inte mer än det .
Det säger jag med eftertryck eftersom jag annars är rädd , och i det avseendet har riktar jag avgörande kritik mot det fleråriga utvecklingsprogrammet , nämligen att det i för liten utsträckning är inriktat på hanteringen av kvoter , att det är ett medel som leder till att särskilt medlemsstater med ett något annorlunda system eller en alldeles utmärkt kontroll över att kvoterna verkligen efterlevs , träffas extra hårt .
I det sammanhanget vill jag yrka starkt för den position fiskeriländerna kring Nordsjön och det nordatlantiska området har .
Herr talman !
Jag håller fast vid att jag hyser stor uppskattning för uppläggningen av Cunhas program , för hans betänkande , men jag har mycket kraftiga principiella invändningar när han lägger fram möjliga sanktioner angående en minskning av kvoterna , även om det bara är tillfälligt .
Det medlet kan inte användas i det här fallet .
Det är en helt annan politik och jag anser att parlamentet principiellt måste förkasta den saken och att vi måste kämpa för att vi i alla fall får en bättre fiskeripolitik med bättre kontroll över vad som händer och sker .
På grundval av detta kan vi också föra en bättre politik .
Det är det första steg som vi måste ta .
Ett andra steg är efterlevandet av kvoterna , det har vi andra medel för .
Det tredje är att ett flerårigt utvecklingsprogram måste vara inriktat på omstrukturering och ingenting annat .
Herr talman !
En särskild gratulation till Cunha för hans utmärkta betänkande .
Kolleger !
Kommissionens rapport går igenom de olika medlemsstaternas arbete och visar att Portugal mycket väl uppfyllt de mål som har fastställts inom samtliga flottsegment , vilket visar en god överensstämmelse mellan informationen i flottregistret och den situation som har presenterats i den portugisiska regeringens rapport .
Angående rapporten om 1997 saknades bara information om fem fartyg i flottan , vilket nu är löst då det bara saknas information om tre fartyg .
Denna aspekt om uppfyllande av målen i de fleråriga utvecklingsprogrammen , som skulle kunna och borde vara positiv , har lett till negativa reaktioner på nationell nivå , dels från fiskerisektorn , dels från pressen och allmänheten generellt sett , eftersom uppfyllandet av målen vanligtvis betyder en minskning av flottans kapacitet och storlek .
Man kan inte straffa dem som uppfyller målen och detta måste förklaras för fiskarna , varför vi föreslår effektiva sanktioner som exempelvis en tillfällig minskning av kvoter för de stater som brutit eller inte uppfyllt de förutsatta fristerna för att lämna in sina uppgifter .
Vi skulle således vilja sätta in sakerna i ett sammanhang : när man säger att vi förstör alltfler fartyg , så stämmer inte det med verkligheten , åtminstone inte om vi jämför med den nuvarande situationen .
I Portugal presenterades , under perioden 1992 till 1995 , 144 nya projekt ; under perioden 1996 till 1999 presenterades 194 projekt , under år 1999 har 40 nya projekt presenterats .
En viktig aspekt som vi dock vill uppmärksamma kommissionen på är följande : omställningen av flottan måste ske med hänsyn till behoven att skydda arbetsvillkoren ombord och de hygienisk-sanitära villkoren för fisken .
Detta kan många gånger kräva ett ökat bruttotonnage .
Slutligen skulle jag vilja be kommissionen , när den fastställer ett eventuell framtida flerårigt utvecklingsprogram V , att inte börja från början utan ta hänsyn till de ansträngningar som redan har gjorts av medlemsstaterna och de resultat som har uppnåtts i tidigare fleråriga utvecklingsprogram .
Herr talman !
Jag vill säga att jag helhjärtat stöder betänkandet som har utarbetats av Cunha .
På samma gång som jag har reservationer , ser jag ingen annan väg framåt .
Det är en intressant tanke att de medlemsstater som har stora flottor i dag byggde upp dessa flottor på femton- och sextonhundratalet .
I Irland känner vi oss djupt förfördelade på grund av storleken på våra kvoter och kapaciteten hos vår flotta .
Vi måste komma ihåg att det när andra sjöfartsnationer - Storbritannien , Spanien , Holland - byggde upp sina flottor på femton- och sextonhundratalet faktiskt fanns en lag som förbjöd fisktransport på irländska skepp .
Så vi gick in i detta århundrade med samma slags båt , den lilla curragh-båten , som St Brendan använde för att segla till Amerika på sjuhundratalet .
Det är därför de fiskare som jag företräder känner sig mycket förfördelade .
Nederländerna har i dag sju gånger så många fartyg över 24 meter som Irland har , även fast vi har mycket större resurser i havet .
Jag vill till protokollet föra det faktum att vi inte är tillfredsställda och säga att vi förmodligen skulle kunna hämta dubbelt så mycket fisk ur de europeiska vattnen jämfört med vad vi hämtar i dag , om vi utnyttjade haven och skyddade och hanterade våra fiskresurser såsom vi borde .
Vi skulle inte få flera arbeten , eftersom vi redan har den kapacitet som behövs , men vi skulle mer än fördubbla de vinster som vi gör för närvarande .
Ett förståndigt system för skydd och återhållsamhet i dag kommer att garantera resurserna för kommande generationer .
När vi har gjort detta och trots det faktum att " relativ stabilitet " har blivit en helig princip här , hoppas jag verkligen att ett land som Irland , vid Atlantens rand , med väldiga resurser , en dag kommer i åtnjutande av en mer rättvisa andel .
Herr talman !
De fleråriga utvecklingsprogrammen för fiskerinäringen har införts för att se till att länder håller sig till överenskomna fångstkvoter .
Eftersom medlemsstaterna inte gjorde det så behövde fiskeflottorna minskas .
I Nederländerna har vi valt en lösning som är typisk för vårt land .
Det har träffats avtal med fiskerisektorn angående en minskning av antalet dagar till havs .
På det sättet behöver inte moderna , lönsamma fartyg tas ur bruk och går företag inte i konkurs och naturligtvis , det allra viktigaste , klarar Nederländerna på det sättet de ålagda fångstkvoterna .
Cunhas betänkande , som jag för övrigt uppskattar , innebär nu att länder som inte håller sig till de fleråriga utvecklingsprogrammen automatiskt måste minska sina fångstkvoter .
Det strider inte endast mot alla rättvisans principer , det är också att spänna hästen bakom vagnen .
Målsättningen med de fleråriga utvecklingsprogrammen är ju att tvinga länder till att fiska inom sina fångstkvoter .
Det vore absurt att ålägga en straffminskning , särskilt en automatisk straffminskning , för ett land som respekterar sina fångstkvoter , som till exempel Nederländerna .
På det sättet kommer medlet att stå över målet .
Det är också för tidigt med en sådan åtgärd .
Nederländerna är ett av de få länder som lämnar tydliga uppgifter om flottkapacitet och fångstkvoter .
Först när det finns ett enhetligt sätt att mäta dessa uppgifter i alla medlemsstater kan man verkligen börja undersöka om alla medlemsstater håller sig till målsättningen .
Avslutningsvis så håller sig Nederländerna samtidigt till arbetstidsdirektivet genom att efterleva fångstkvoterna genom att minska antalet dagar som båtarna ligger ute .
Även om fiskerisektorn egentligen inte omfattas av det direktivet så har naturligtvis även fiskare rätt till en lämplig vilotid .
En minskning av antalet dagar till havs kan bidra till det .
Herr ordförande !
Min delegation skall rösta mot betänkandet om punkt 6 i resolutionen antas . .
Herr talman !
Först och främst vill jag tacka Cunha för ett utmärkt betänkande och gratulera mig själv till resolutionen om kommissionens årsrapport om det fleråriga utvecklingsprogrammet .
Jag vill påpeka att såväl detta betänkande som tidigare av Cunha utarbetade resolutioner med anledning av den bristande fullgörelsen av de fleråriga programmen har varit kommissionen till stor nytta vid utformningen av nya lagar , särskilt inför tillämpningen av FIUF-fonderna som godkänts för nästkommande år .
Kommissionen håller helt och hållet med Cunha och andra talare i att de fleråriga utvecklingsprogrammen är av stor vikt för att kunna säkerställa framtiden för gemenskapens fiskeflotta .
Vissa punkter vill jag dock poängtera .
För det första hur mätning skall utföras - en nyckelfråga när det gäller hur de olika länderna verkligen följer FUP - även om det är riktigt att man ännu inte har lyckats uppnå en fullständig harmonisering av mätenheterna vid övergången från ett system till ett annat , så håller kommissionen på med detta och vissa initiativ har tagits .
Bland annat har man beställt en uttömmande rapport i ämnet från en extern expert , Seafish Industries Authorities , som har besökt behöriga myndigheter i de olika länderna för att på lämpligt sätt studera hur mätningarna skall harmoniseras .
Genom att basera sig på detta betänkande tillsammans med de rapporter och arbeten som utformats av gemenskapsinspektörerna så kommer kommissionen att utarbeta ett förslag till revision av mätningsförordningen , det vill säga ett revisionsförslag för övergången mellan FUP III och FUP IV .
Ärade kollegor , herr talman , jag vill också tillägga att kommissionen samarbetar med Europeiska standardiseringsorganisationen ( CEN ) för att fastställa en gemensam standard för mätning av drivkraft , ett annat sätt att mäta varje flottas fiskekapacitet .
När vi vet hur vi bättre skall definiera FUP och när vi vet hur varje flottas fiskekapacitet skall mätas så kommer vi till den mest polemiska frågan .
Kontrollen av hur de fleråriga utvecklingsprogrammen följs , den kontroll som rådet fastställer efter kommissionens förslag .
Kommissionen är inte nöjd med hur den här frågan handläggs , och även om vissa framsteg gjorts så har man inte gjort allt det som kommissionen föreslagit .
Framsteg har gjorts i och med att de offentliga stöden har tagits bort vilket är ett effektivt instrument , åtminstone för en del medlemsstater som har ändrat hållning och börjat tillhandahålla mera information .
Effektivare fleråriga utvecklingsprogram har tagits fram och därför kan man säga att framsteg gjorts .
Den nya strukturella politiken inom fiskerisektorn för perioden 2000-2006 inkluderar helt klart nya bestämmelser beträffande påföljder som - en gång för alla - skall ge kommissionen medel för att av medlemsländerna lättare kunna kräva fullgörelse av de olika FUP .
Låt mig påpeka för er som ansåg att de godkända sanktionerna var otillräckliga att detta inte berodde på kommissionen .
Kommissionen hade föreslagit kompletterande påföljder men detta avslogs av rådet .
Tilläggssanktioner som till exempel att länder som inte på ett ändamålsenligt sätt följer FUP skulle förhindras att delta i nya fisketurer i tredje land finansierade av gemenskapsfonderna .
En sådan åtgärd hade varit mycket effektiv men den avslogs av rådet .
Det är med andra ord inte kommissionen som inte vill använda sig av effektivare metoder för att nå bättre fullgörelse .
Det är rådet .
Kommissionen är beredd att gå vidare och vad som saknas är att rådet visar en liknande vilja .
Med anledning av polemiken kring artikel 6 , måste jag säga att vissa problem av juridisk karaktär uppstår .
Eftersom det bara är fråga om en temporär reträtt så skulle man kunna ta något sådant i beaktande .
Det finns dock andra system men rådet vill inte godkänna dessa heller .
Vi tvivlar på att rådet kommer att ändra sig och godta ett sådant förslag .
Ändrar de inställning kommer dessa eller andra förslag att välkomnas .
Andra förslag kommer nog att läggas fram eftersom kommissionen redan har gjort sitt och det var rådet som satte sig på tvären .
Ärade kollegor , vi måste förvisso komma ihåg att det till syvende och sist ofta är producenterna som bestraffas .
Om vi drar en parallell mellan jordbruk och fiske - vilket vi mycket väl kan göra - så kommer en viss typ av sanktioner att beröra jordbrukaren , som plötsligt får se sin inkomstkälla minskas .
En minskning av flottan i ett land innebär givetvis en uppoffring för den befolkning som lever vid och av havet och som berörs av en sådan minskning .
Vissa åtgärder berör den sociala sektorn och varje land - samt gemenskapen - måste vidta kompletterande åtgärder för att mildra effekterna .
Ärade kollegor , det är med fullgörelsen av FUP , särskilt när det gäller fiskekvoter och en rationell hantering av fiskeresurser , som vi verkligen sätter den europeiska fiskerisektorns framtid på spel .
Jag tackar och lyckönskar än en gång Cunha för betänkandet , och jag upprepar att när det gäller fullgörelse och sanktioner så är det kommissionen som har lagt fram positiva förslag och andra som inte har velat ha dem och att kommissionen givetvis kommer att fortsätta att försöka se till att medlemsländerna bättre uppfyller sina åtaganden .
Tack , kommissionär Palacio !
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i dag kl .
12.00 .
 
Energieffektivitetskrav för förkopplingsdon till lysrör Nästa punkt på föredragningslistan är debatt om betänkande ( A5-0102 / 1999 ) av Turmes för utskottet för industrifrågor , utrikeshandel , forskning och energi om förslaget till Europaparlamentets och rådets direktiv om energieffektivitetskrav för förkopplingsdon till lysrör ( KOM ( 1999 ) 296 - C5-0010 / 1999 - 1999 / 0127 ( COD ) ) . .
( DE ) Herr talman , fru kommissionär , ärade kolleger !
Varför ett europeiskt direktiv om effektiviteten i lysrör ?
Vi använder årligen 130 miljoner sådana lysrör i de 15 EU-länderna , i synnerhet i kontorsbyggnaderna , där två tredjedelar av ljuset numera kommer från lysrör .
1992 genomförde Europeiska kommissionen med anledning av konferensen i Rio en undersökning om vilka konkreta åtgärder man i våra länder kan vidta för att skydda klimatet .
Då upptäcktes att en av least-cost-åtgärderna inom EU skulle vara effektivare lysrör .
Man skall vara medveten om att dessa lampor lyser tio timmar per dag , fem till sju dagar i veckan , 50 veckor per år och under många år och att även en mycket liten effektivitetsskillnad - om den så bara är på tre eller fem watt - under årens lopp gör väldigt mycket för elförbrukningen .
Kommissionen inledde 1993 förhandlingar med CELMA , sammanslutningen för belysningstillverkare , och genomförde 1996 en studie för att skapa en vetenskaplig bas för ett beslut .
I denna studie från 1996 kalkyleras det med ett flertal scenarier , och det mest långtgående scenariot , enligt vilket alla magnetiska förkopplingsdon så småningom helt försvinner från marknaden och the best available technology , de elektroniska förkopplingsdon som i dag innehar 20 procent av marknaden , dominerar hela marknaden , skulle innebära 250 terawattimmar , 250 miljarder kilowattimmar för det sammantagna EU-området .
Jag kommer från Luxemburg .
Luxemburgs totala elförbrukning - för industri , hushåll , kontorsbyggnader - uppgår till 6 terawattimmar per år .
Med hjälp av direktivet skulle vi alltså årligen kunna spara dubbelt så mycket som Luxemburgs totala elförbrukning , dvs. det är inte så irrelevant som det kan tyckas vid en första anblick .
Kommissionen lade 1999 fram en proposition .
I förslaget lägger man sig rentav under minimiscenariot i studien som kommissionen själv gav i uppdrag 1996 .
Detta beror på att phasing out-momentet inte genomförs konsekvent för alla magnetiska förkopplingsdon och att olika magnetiska don därmed skulle bli kvar på marknaden , och att vi sparar in 100 miljarder kilowattimmar mindre under de kommande åren .
Därför bör vi som parlament förbättra kommissionens proposition .
Det finns ekologiska argument , vilka jag redan har åberopat .
Det finns dock även ett tekniskt , finansiellt argument .
Industrin själv har på grundval av det aktuella lagförslaget från kommissionen försökt uppskatta vilka investeringssignaler som ges till marknaden för förkopplingsdon och slagit fast att 50 procent av förkopplingsdonen om 5-8 år därmed skulle komma från de bästa magnetiska förkopplingsdonen , dvs. att vi egentligen ger en felaktig signal till marknaden .
I stället för att styra in hela investeringsvolymen på the best available technology , de elektroniska förkopplingsdonen , skulle en stor del av investeringarna gälla den näst bästa tekniken .
Man kan således föreställa sig att industrin , ifall man under de kommande 3-4 åren investerar i den näst bästa tekniken , om 5-6 år - då vi är på gång med en review - kommer att värja sig ännu mycket starkare än i dag mot att häva just dessa nyinvesteringar .
Och nu litet background för det internationella sammanhangets skull : I USA räknar man med en phase out av alla magnetiska förkopplingsdon fram till år 2010 .
Vårt förslag - och här vill jag tacka skuggföredragandena från de andra partierna , McNally , Rovsing och Beysen - skulle inte innebära något annat än vad som redan är på gång i USA .
Herr talman !
Jag tackar föredraganden för upplägget , vilket jag fullständigt stöder .
Jag tackar för ett gott samarbete mellan grupperna , genom vilket vi nått fram till kompromisser som jag tycker är ansvariga , korrekta och lämpliga .
Vi står därför bakom dem i vår grupp .
Varför befattar vi oss med detta ?
Ja , för att säga det mycket kortfattat handlar det alltså om att begränsa det utsläpp av koldioxid som härrör från människors handlingar .
Vi vet att efterhand som man får en högre levnadsstandard i Asien , kommer 1,4 miljarder kineser och 1 miljard indier att börja använda mer och mer energi och detta betyder att deras energiförbrukning från nuvarande 10 procent av EU : s genomsnittliga energiförbrukning kommer att öka våldsamt , när de efterfrågar vanliga , grundläggande bekvämligheter som t.ex. varmvatten och kanske också luftkonditionering , transporter och en modern industri .
I Rio åtog vi oss att skydda klimatet .
Genom detta dokument uppfylls detta syfte till fullo .
Vi kan se att av den koldioxid som härrör från människors handlingar , kommer 30 procent från elproduktionen .
Och 35 procent av all energianvändning i EU kommer från elektricitet .
De långa , raka lysrören står i EU för 53 procent av elförbrukningen till belysning .
Och om vi lyckas genomföra det enligt planering , kommer vi år 2020 att spara 6 miljoner ton koldioxidutsläpp per år .
Vi kommer att spara 10 procent av elförbrukningen till lysrörsbelysning , och i pengar räknat blir det en besparing på 250 miljoner euro per år .
Detta förslag kan alltså få ganska avsevärda effekter på klimatet och på ekonomin och genom att vi genomför det enligt förslaget , ger vi vår industri lång tid att ställa om sig .
Turmes tog upp detta och jag kan påminna mig om att i varje fall sedan 1992 har industrin känt till att runt år 2009 kommer magnetiska förkopplingsdon mer eller mindre att vara förbjudna .
Så det är inget nytt i det vi genomför .
I den kompromiss vi har utarbetat har vi varit överens om att genomföra en effektivisering .
Vår vilja har varit att skydda klimatet .
Vi har velat erhålla ekonomiska fördelar och vi har velat se till att det gradvisa borttagandet som sker inte belastar vanliga konsumenter i vanliga hem onödigt mycket vad gäller investeringar , som inte kan återbetalas , samtidigt har vi sett till att vi i den nordliga delen av unionen , i norra Finland , i norra Sverige , i norra Norge , på Grönland och andra platser där elektroniska förkopplingsdon inte fungerar , kan fortsätta att använda magnetiska förkopplingsdon .
I det stora hela är det ett lysande förslag och jag rekommenderar att vi allihop ställer oss bakom det , just som avtalats i grupperna , och stöder det .
Herr talman !
Det gläder mig att ni finner denna debatt bildande och upplysande .
Debatterna är inte alltid spännande ; det är mycket intressantare att tala om dramatiska väderförhållanden och stormar i Frankrike .
Men om vi vill få ett slut på sådana händelser , är det den här sortens detaljerat , tekniskt arbete som vi måste uträtta .
Jag skulle vilja gratulera Turmes för hans mycket grundliga arbete , hans tekniska sakkunnighet och hans beredvillighet att delta i särskilda kompromissdiskussioner med ledamöter från andra grupper .
Det uppskattas , och jag anser att det är på ett sådant ansvarsfullt sätt som vi bör arbeta här i parlamentet .
Om vi tar våra Kyotoåtaganden och andra åtaganden på allvar och om vill förhindra tragiska väderhändelser , måste vi arbeta med åtminstone det ena ögat på klockan .
Det är åtta år sedan förhandlingar inleddes , med den berörda industrin och med energiexperter , om hur vi skulle kunna använda belysningssektorn för att spara elektricitet .
Det finns många skäl att göra det - det är en extremt förståndig investering för företagen i Europeiska unionen att ha en energieffektiv belysning .
Vi måste ha en inre marknad utan omotiverade , hindrande handelsbarriärer .
Våra företag runtom den inre marknaden måste arbeta på samma villkor ; vi måste ha den berömda jämna spelplanen som mål och alltid ta hänsyn till särskilda nationella intressen och förhållanden .
Elektricitet , påminner oss kommissionen om , står för 35 procent av vår totala förbrukning av primärenergi och är upphov till 30 procent av de koldioxidutsläpp som orsakas av människan .
Att ta itu med denna sektor , liksom med transportsektorn , är av största vikt .
Det är därför lämpligt att vi undersöker miniminormer för effektivitet på varje område där energi förbrukas .
Vi har med framgång undersökt hushållskokare och kokare för industrin , kylskåp och frysar , och vi har ett antal frivilliga överenskommelser - som jag möjligen har reservationer om - på andra sektorer för hushållsapparater .
Om jag får citera från en undersökning som har genomförts i Storbritannien , vid vårt mycket välkända centrum för byggnadsforskning : " Att utarbeta prestandanormer , särskilt för förkopplingsdon till lysrör , ter sig enligt denna undersökning vara en av de mest effektiva åtgärder som EG kan vidta för att minska energiförbrukningen för belysning i byggnader för kommersiella ändamål , och det är följaktligen värt ytterligare övervägande och utveckling . "
Detta mycket högt ansedda forskningscentrum beslutade att detta var en sektor som vi borde arbeta med .
Ett problem är att de som köper lysrör inte nödvändigtvis är samma personer som använder dem .
De som investerar i byggnader är inte samma personer som kommer att betala elräkningarna i framtiden .
Det väldiga antalet lysrör medför emellertid att vi måste se till att dessa köpare måste göra förnuftiga köp , genom att se till att produkterna på marknaden uppfyller högsta möjliga normer .
Vi talar enbart om nyproducerade förkopplingsdon till lysrör .
Vi föreslår inte att vartenda ett måste ersättas i morgon eller nästa vecka .
Det skulle vara ett absurt sätt att gå framåt .
Vi föreslår att de nuvarande lysrören , allt eftersom de tar slut och ersätts under de närmaste 15-20 åren , på ett mycket gradvis , väl avvägt och välövervägt sätt ersätts med den bästa möjliga tekniken .
En mycket lång anpassningsperiod , det är så vi arbetar i Europeiska unionen .
Vi hoppar inte på våra företag med överraskningspaket som de inte har förvarnats om och som skulle orsaka dem ansenliga svårigheter .
Turmes har verkligen varit resonlig .
De 800 personer som är sysselsatta med tillverkningen av magnetiska förkopplingsdon kommer inte att bli av med jobben i nästa vecka .
Det kommer att finnas gott om tid för en infasningsperiod .
Vi i den socialistiska gruppen är emot de extra ändringsförslag som har lagts fram .
De ligger inte i linje med målen i betänkandet .
Men vi stöder de ändringsförslag som vi undertecknade som en del av kompromissen , av vilka många - och jag är säker på att kommissionen skulle hålla med om det - lägger till förnuftiga definitioner .
Jag hoppas att kommissionären kommer att tala om för oss att detta bara är en del i hennes målsättning att öka energieffektiviteten inom Europeiska unionen och göra våra löften till mer än politiska rubriker .
Herr talman , fru kommissionär , kolleger !
Det här betänkandet , som Turmes arbetat fram med stor noggrannhet , verkar vid första anblicken vara en teknisk angelägenhet .
Ändå har det här betänkandet , så vitt jag kan se , mycket större konsekvenser , vilket redan understrukits av kollegerna .
Å ena sidan är det det första betänkande detta årtusende som kommer att bidra till en sparsammare energiförbrukning , och ingen skall ifrågasätta att överlevnadschanserna för vår planet i det här nya årtusendet i hög grad kommer att avgöras av på vilket sätt vi kommer att använda energin i framtiden .
Av den anledningen får man inte aningslöst förbigå det här initiativet .
Å andra sidan anser jag att det sätt på vilket det här betänkandet arbetats fram , via förhandlingar med den berörda industrin och med politiker och med kommissionen , är ett bra exempel på vad man på franska skulle kalla " cohabitation " .
Därmed menar jag att de rådfrågningar och rundabordssamtal som föregick förslaget till direktiv har lett till enighet mellan näringslivet och kommissionen .
Betänkandet är , i föreliggande form , även resultatet av kompromissändringsförslag som godkänts av de viktigaste politiska grupperna och jag ansluter mig till det som den föregående talaren , McNally , sade om att det är ett sätt att arbeta som borde få mer utrymme i framtiden .
I kompromissändringsförslagen anges särskilt långa övergångsperioder .
Det innebär i princip att näringslivet i praktiken får tio år på sig för att genomföra alla de anpassningar som behövs .
Dessutom bör tilläggas att man från näringslivets sida redan sedan år 1992 visste att förändringarna var oundvikliga .
Dessutom är det också bra att veta att de magnetiska förkopplingsdonen definitivt måste vara utbytta först från och med år 2009 .
Betydelsen av det här betänkandet , herr talman , ligger samtidigt i den viktiga effekt som det här direktivet har för sysselsättningen för tusentals arbetstagare samt även i uppmärksamheten för störningen av konkurrenspolitiken .
Om övergångsperioderna skulle göras för korta så är det ju klart att inte endast en fullständig produktionslinje utan även producenten skulle hamna i farozonen eftersom den senare inte skulle ha någon möjlighet att i tid anpassa produktionslinjen .
Det skall självklart vara så att förhandlingar hålls regelbundet under genomförandet av direktivet , så att de som hittills inte varit positivt inställda till bytet av förkopplingsdon får möjlighet att förstå utvecklingsprocessen .
Genom att göra en avvägning mellan de olika intressena och genom ett nära samarbete med de olika intressenterna har parlamentet lyckats lägga fram ett tydligt och väl underbyggt lagstiftningsarbete .
Mina gratulationer till kollega Turmes för det .
Herr talman !
Det här betänkandet handlar om en mycket teknisk fråga , men det är av stor betydelse såväl för sparandet av energi som för den europeiska sysselsättningen .
Föredraganden har gjort ett utmärkt arbete för att klargöra betänkandets energieffekter , men samtidigt har man inte i tillräcklig utsträckning beaktat att genomförandet av betänkandet skulle skapa arbetslöshet i Europa , mest i Tyskland , men också i Finland , Österrike , Italien och Spanien .
I lysrör används två typer av förkopplingsdon som påverkar energins effektivitet .
Magnetiska förkopplingsdon alstrar mycket ljus och mycket värme .
I nordliga länder sparar denna värme uppvärmningsenergi och är inte enbart spillvärme .
Elektroniska förkopplingsdon producerar bättre ljus och mindre värme och är vad gäller energins effektivitet klart bättre än de magnetiska förkopplingsdonen .
Framtiden är deras om de kan göras lika konkurrenskraftiga ekonomiskt som de magnetiska förkopplingsdonen .
Företaget Philips har säkert gjort rätt i att investera i den här tekniken .
Dess produkter borde dock inte genom politiska tvångsåtgärder göras till enda europeisk standard .
Tvärtemot kommissionen och rådet föreslår Turmes att de magnetiska förkopplingsdonen till lysrör skall förbjudas .
Om betänkandet godkändes skulle parlamentets ståndpunkt utplåna den europeiska industrin på området .
I resten av världen skulle man nog fortsätta att tillverka och använda magnetiska förkopplingsdon , som är nödvändiga under sådana klimatförhållanden som jag kommer ifrån : Där det är kallt eller fuktigt kan man bara använda magnetiska förkopplingsdon .
På grund av förbudet skulle produktionen av magnetiska förkopplingsdon flyttas från Europa till utvecklingsländerna .
I USA har man redan erfarenheter av detta .
Vill man behålla arbetstillfällen i Europa kan man inte godkänna Turmes betänkande med avseende på de delar som kollegan Westendorp y Cabezas ändringsförslag behandlar .
Jämfört med magnetiska förkopplingsdon är produktionskostnaderna för elektroniska förkopplingsdon tio gånger så stora , och skonandet av naturen skall också ses ur materialförbrukningens och återvinningens synvinkel .
Herr talman , jag uttalar mig för TDI-gruppen även om jag talar på en av dess beståndsdelars vägnar .
Vi har tillfrågats om problemet med förkopplingsdon till lysrör .
Vad handlar det om ?
Elströmmen i lysrör såsom de som belyser oss där uppe ovanför våra huvuden , regleras och stabiliseras av små apparater som kallas för förkopplingsdon .
Dessa förkopplingsdon tillverkas sedan femtio år tillbaka av en kopparrulle i en plåtdosa .
De kallas " ferromagnetiska " .
Men det finns nu elektroniska förkopplingsdon .
Det sägs att de traditionella ferromagnetiska donen medför en energiförlust , i synnerhet genom ett motståndsfenomen .
Förlusten sägs vara ända till 8 watt per timme medan de elektroniska donen bara förlorar 3 watt .
Med dem kan således en besparing på 5 watt göras , säger man , och genom att multiplicera med 130 miljoner förkopplingsdon sparas miljoner ton energi , det blir mindre koldioxid , mindre växthuseffekt och mänskligheten andas bättre .
Vi måste därmed på åtta år överge de ferromagnetiska förkopplingsdonen för elektroniska .
Turmes säger tyvärr inte till oss att de elektroniska förkopplingsdonen har kortare livslängd än de ferromagnetiska .
Vi måste således tillverka fler med mer energi som går åt och besparingarna nyss försvinner delvis .
De elektroniska förkopplingsdonen tillverkas dessutom med transistorer som innehåller tunga metaller , såsom tantal , germanium och till och med arsenik för att inte tala om plast , dvs. icke biologiskt nedbrytbara förorenande ämnen , medan koppar och plåt från de magnetiska donen är biologiskt nedbrytbara .
Med andra ord , för att göra en mindre uppenbar energibesparing än till synes slänger våra gröna kolleger ut tunga metaller och arsenik i naturen .
Förutom att man ökar föroreningarna ökar man för övrigt på samma gång arbetslösheten eftersom de komponenter som ingår i elektroniktillverkningen och de maskiner som tillverkar dem inte är europeiska .
Följaktligen för att undvika importkostnader skall våra industrier omlokalisera sig och således minska arbetstillfällena .
Genom att försiktigt vilja spara energi med elektronik medan våra industrier bara begär ett gradvist och selektivt förbud , får vi sammanlagt i bästa fall en besparing men med utsläpp av förorenande ämnen och arbetslöshet i tillägg .
Och man tar inte itu med den verkliga frågan om slöseri , det vill säga glödlampor som förlorar upp till 50 watt jämfört med lysrör .
Men glödlampor tillverkas ju av två multinationella företag , Philips och Osram .
Och kanske det blir kontakt mellan Europeiska kommissionens anhängare av globalisering , det dunkla gröna multinationella partiets anhängare av globalisering och de gränsöverskridande industriföretagen , men jag begär inte att man belyser frågan fullt ut .
Herr talman , mina damer och herrar !
Jag blickar uppåt här i salen och kan konstatera att vi är omgivna av väldigt många förkopplingsdon .
Jag tror att denna sal är en förebild för hur neonrör och förkopplingsdon samarbetar .
Jag är säker på att vi redan har de energisnåla elektroniska lamporna här , för det har ju bevisats att de elektroniska förkopplingsdonen betalar sig inom ett eller ett par år .
Vi har alltså ett mycket bra return on investment , och därför går egentligen alla moderna byggare och planerare redan nu över till de elektroniska förkopplingsdonen .
Det förhåller sig för närvarande så att marknaden inte alls klarar av att producera så många apparater som egentligen skulle behövas .
Det egentliga problemet ligger i att tekniken är så modern och så attraktiv att industrin faktiskt inte kan framställa erforderliga mängder för den närmaste tiden .
Detta är naturligtvis också ett problem , att vi måste träffa en överenskommelse för att instrumenten skall finnas tillgängliga i tid , eftersom vi annars kommer att stå där med en viss brist .
Om det inte längre går att tillverka de magnetiska donen och de elektroniska samtidigt inte finns i tillräckligt antal kan det uppstå problem på marknaden .
Men jag är ändå för en legislativ reglering , även om jag länge har funderat kring huruvida det alls är meningsfullt med ett europeiskt direktiv för förkopplingsdon .
Jag är för detta eftersom jag anser att vi framdeles bör satsa på mer forskning i tekniken i fråga .
Vi bör arbeta för att garantera att investeringarna också i framtiden skall gälla de elektroniska donen .
Redan nu är detta en självklarhet för marknaden .
Men jag tror absolut att direktivet kan vara en sporre till att investera ännu mer och ännu snabbare och därmed till att tjäna stora pengar .
Herr talman !
De talare som redan har yttrat sig visade verkligen att de är kompetenta när det gäller ett ämne som är så extremt tekniskt som förkopplingsdon till lysrör .
Men det verkar som om debatten inte har haft så stor intresse och jag frågar mig hur många av mina kolleger som faktiskt kan rösta med sakkunskap i frågan , med tanke på att när det gäller en persons allmänbildning - de kunskaper man får genom studier , genom privata erfarenheter eller genom de politiska erfarenheter man gör som parlamentariker - så är det inte ofta man hittar djupgående kunskaper när det gäller förkopplingsdon till lysrör .
Jag frågar mig därför om den här typen av frågor måste debatteras i kammaren eller om det kanske inte hade varit bättre att bara hänvisa till de regler som finns och diskutera frågorna i utskottet .
Vissa frågors extremt tekniska natur gör det i själva verket omöjligt att rösta på ett kunnigt sätt om man nu inte skall gå efter de vanliga kryssen och strecken på listor som utarbetats av någon annan .
Men detta är att förringa parlamentarikernas verksamhet !
Man undrar dessutom om det verkligen är nödvändigt att parlamentet sysslar med så här komplicerade och extremt tekniska frågor eller om det inte i stället skulle vara bättre , vilket sker i de olika nationella lagstiftningarna , att ge andra organ behörighet att besluta i dessa frågor , med tanke på att de politiska återverkningarna - detta har vi fått höra även av de talare som redan har yttrat sig - är minimala .
Låt mig också göra ett påpekande när det gäller den så kallade rena energin , något som verkar ha undgått många talare .
Det är inte sant att elenergin är en ren energi .
Det är klart att om jag värmer upp mitt hus med elradiatorer i stället för vattenfyllda element som värms med olja , så blir föroreningarna mindre i städerna , men om man tänker på , vilket också påpekas i betänkandet , att för att producera elenergi så släpper vi i atmosfären ut 30 procent av all koldioxid , så är det kanske dags att även den allmänna opinionen omvärderar sina kunskaper och sina övertygelser och , framför allt , att medierna blir tydligare när ett gäller vilka energiformer som verkligen är rena och vilka som i stället inte är det .
Herr talman !
Först och främst vill jag lyckönska föredragande Turmes för ett utmärkt betänkande samtidigt som jag vill tacka alla talare och parlamentet för det stöd som givits förslaget , ett förslag som kommissionen tror i hög grad kommer att bidra till ökad energieffektivitet där målet är att spara 20 procent av elförbrukningen för den tredje sektorn .
För att substantiellt förbättra effektiviteten hos slutanvändaren är detta nödvändigt och därmed bidrar vi till att fullfölja våra åtaganden från Kyoto .
I förslaget har man antagit ett omsorgsfullt utarbetat projekt för att förbättra effektiviteten utan att detta medför en outhärdlig överbelastning för tillverkarna av förkopplingsdon .
Jag vill nämna , ärade kollegor , att precis som en av talarna sade så har vi innan förslaget godkändes rådfrågat och talat med den berörda sektorn .
Ärade kollegor , vi utgår från ett förslag i olika steg .
Den första nivån som tas i bruk ett år efter direktivets antagande innebär en progressiv minskning av förkopplingsdon med låg effektivitet .
Därefter övergår vi till nivå två som är mera krävande och där konventionella förkopplingsdon progressivt minskas och bruket av högeffektiva förkopplingsdon blir obligatoriskt .
För att ni skall förstå vad detta innebär måste jag säga att dagens konventionella förkopplingsdon står för cirka två tredjedelar av den totala försäljningen , vilket medför att den andra nivån kommer att få mycket stora effekter och otvivelaktigt återverka på industrin och att vi därför föreslår en övergångsperiod på fyra år .
När det gäller de ändringsförslag som lagts fram så gläder det mig , ärade kollegor , att få tala om att kommissionen kan godkänna alla som lagts fram av utskottet för industrifrågor , utrikeshandel , forskning och energi , förutom ändringsförslag 1 , 17 , 19 och 20 om införandet av en tredje automatisk effektivitetsnivå .
Kommissionen håller med om att det krävs en dynamisk framställning och därför förutser man i förslaget en eventuell tredje fas .
Vi menar dock att det just nu är svårt att bestämma hur en sådan tredje fas skall se ut .
Vi menar att det är bättre att utvärdera den tekniska och ekonomiska situationen när den andra fasen träder i kraft och då bestämma , genom att rådfråga berörda parter , om fas tre skall genomföras , hur den skall genomföras , vilka de tekniska definitionerna är samt vilka krav som skall ställas och när den skall sättas i gång .
Kommissionen kan följaktligen även godkänna andra delen av ändringsförslag 23 , men inte den första delen .
På samma sätt kan kommissionen godkänna första delen av ändringsförslag 1 , i en annorlunda tappning .
Vi är dessutom eniga vad gäller ändringsförslag 12 så att medlemsländerna på ett effektivt sätt kan tillämpa det .
De ändringsförslag som syftar till att klargöra att alla förkopplingsdon som marknadsförs som fristående komponenter eller inmonterade i lysrör är täckta av förslaget , det vill säga ändringsförslag 3 , 4 , 5 , 6 , 7 , 8 , 9 , 10 , 11 , 13 , 14 , 21 och 22 , och som jag redan nämnt godkänner kommissionen alla .
Ändringsförslag 2 godkänns också eftersom kommissionen håller med om att den typen av förkopplingsdon skall uteslutas .
Ändringsförslag 15 och 16 där övergångsperioden förlängs till 18 månader godkänns också .
Avslutningsvis godkänner kommissionen ändringsförslag 8 om hur effektivitetsnormerna vid internationella forum skall marknadsföras .
Herr talman , ärade kollegor , jag har sammanfattat kommissionens ståndpunkt .
Jag tackar än en gång föredragande Turmes som har genomfört ett utmärkt arbete och jag förlitar mig på att rådet kan anta en gemensam ståndpunkt som snabbt kan lösa den här frågan .
( Applåder ) Tack , fru de Palacio !
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i dag kl .
12.00 .
 
OMRÖSTNING Herr talman !
En ordningsfråga .
Den har att göra med mitt betänkande om kvinnor och vetenskap .
Debatten kan äga rum i kväll , men det kommer inte att vara möjligt att rösta om betänkandet i morgon , på grund av extremt allvarliga och vilseledande översättningsmisstag , framför allt i den franska versionen .
Jag skulle vilja be er att klargöra att så snart en rättad version av ändringsförslagen och mitt betänkande finns tillgängliga , kommer omröstningen att äga rum under den närmast följande sammanträdesperioden .
Det är tyvärr inte möjligt att genomföra omröstningen i morgon , eftersom översättningen , särskilt till franska , har så väldigt stora brister .
Låt mig då bara bekräfta detta .
Debatten om McNallys betänkande kommer att äga rum i kväll , men omröstningen kommer inte att äga rum förrän under den korta sammanträdesperioden i Bryssel .
Betänkande ( A5-0102 / 1999 ) av Turmes för utskottet för industrifrågor , utrikeshandel , forskning och energi om förslaget till Europaparlamentets och rådets direktiv om energieffektivitetskrav för förkopplingsdon till lysrör ( KOM ( 1999 ) 296 - C5-0010 / 1999 - 1999 / 0127 ( COD ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Gemensamt resolutionsförslag om oljeutsläpp i Frankrike ( Parlamentet antog den gemensamma resolutionen . )
Gemensamt resolutionsförslag om stormar i Europa ( Parlamentet antog den gemensamma resolutionen . )
Gemensamt resolutionsförslag om fredsprocessen i Mellanöstern Före omröstningen : Herr talman !
Det här ändringsförslaget gäller endast ett misstag som smugit sig in i resolutionstexten , punkt 5 .
Med mitt ändringsförslag vill jag återställa den text som vi hade kommit överens om vid utarbetandet av den gemensamma resolutionen .
Det gäller alltså ett misstag som vi försöker rätta till med det här ändringsförslaget .
Herr talman !
Jag beklagar att jag nu gör något som jag normalt inte brukar göra , nämligen ta till orda om ändringsförslag .
Kollegan de Clercq har satt stenen i rullning .
Därmed blir jag tvungen att ta ställning .
Vi har avtalat texten så som den nu står i tryck .
Det gäller vår uppmaning till Israel att lämna de ockuperade områdena i Libanon .
Enligt avtalet skulle texten se ut som den nu föreligger .
Nu vill liberalerna och kanske även andra här i salen stryka den mening som innehåller uppmaningen till Israel om att dra sig tillbaka från Libanon .
Det är deras fulla rätt att göra så , men vi kan inte påstå att vi har avtalat något sådant .
Vi har avtalat det som står i texten .
Som ni helt korrekt säger , debatterar vi inte ändringsförslagen .
Så låt oss nu fortsätta omröstningen .
( Parlamentet antog den gemensamma resolutionen . )
Gemensamt resolutionsförslag om internationella kapitalflöden ( Parlamentet förkastade det gemensamma resolutionsförslaget . )
Resolutionsförslag ( B5-0089 / 2000 ) av Wurtz m.fl. för GUE / NGL-gruppen om beskattning av kapitalbetalningar ( Parlamentet förkastade resolutionsförslaget . )
Resolutionsförslag ( B5-0090 / 2000 ) av Goebbels m.fl. för PSE-gruppen om införandet av en skatt på kapital ( " Tobinskatt " ) ( Parlamentet förkastade resolutionsförslaget . )
Resolutionsförslag ( B5-0091 / 2000 ) av Jonckheer m.fl. för Verts / ALE-gruppen om kapitalskatt ( Tobinskatt ) ( Parlamentet förkastade resolutionsförslaget . )
Resolutionsförslag ( B5-0092 / 2000 ) av Cox m.fl. för ELDR-gruppen om Tobinskatten ( Parlamentet förkastade resolutionsförslaget . )
Betänkande ( A5-0096 / 1999 ) av Cunha för fiskeriutskottet om den årliga rapporten till rådet och Europaparlamentet om resultatet av de fleråriga utvecklingsprogrammen för fiskeflottorna vid utgången av 1997 ( KOM ( 1999 ) 175 - C5-0109 / 1999 - 1999 / 2112 ( COS ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Röstförklaringar Betänkande ( A5-0102 / 1999 ) av Turmes Herr talman !
Som företrädare för Pensionärspartiet röstade jag för energisparåtgärderna som rör förkopplingsdon till lysrör , även om jag röstade för ett antal ändringsförslag som emellertid inte antogs av parlamentet .
Jag håller med om att vi skall spara energi - i själva verket läser jag sedan en tid tillbaka de betänkanden som skall diskuteras i parlamentet i ljuset från ett stearinljus för att kunna ge mitt blygsamma bidrag till energisparandet - jag anser att vi naturligtvis skall spara energi , men jag anser också att vi måste vara förnuftiga nog att förstå att detta inte får leda till att vi totalt avskaffar alla de verksamheter som ger de europeiska medborgarna sysselsättning . .
( FR ) Kommissionens förslag till direktiv om förkopplingsdon till lysrör syftar till att förbättra deras effektivitet och att minska energiförbrukningen .
I det föreslås att åtgärder vidtas gradvis och balanserat .
Genom att godkänna flera ändringsförslag respekterar inte utskottet för industrifrågor , utrikeshandel , forskning och energi denna balans eftersom det vill avskaffa tillverkning och saluföring av ferromagnetiska förkopplingsdon endast till fördel för elektroniska förkopplingsdon .
Detta maximalistiska tillvägagångssätt tar inte hänsyn till samtliga tekniska och vetenskapliga argument såväl på energibesparingsnivå som i fråga om tekniska framsteg .
Den verkar , till exempel , vara ovetande om att det finns ferromagnetiska förkopplingsdon med låg energiförbrukning som har sin fulla plats på marknaden .
Vad som är ännu allvarligare är att utskottet för industrifrågor , utrikeshandel , forskning och energi är fullständigt ovetande om förslagets återverkningar på sysselsättningen .
Att upphöra med tillverkning av ferromagnetiska förkopplingsdon riskerar att medföra stängning av många produktionsenheter och många permitteringar , liksom , till exempel , i fabriken Vossloh-Schwabe i Colmar .
Därför röstade jag emot det slutliga betänkandet efter godkännandet av många ändringsförslag som skulle vara mycket farligt för sysselsättningen inom sektorn om de tillämpades .
Jag vill uppmana rådet att förkasta de ändringsförslag som just godkänts .
Gemensam resolution om oljeutsläpp i Frankrike De franska västliga kustområdena är nu nedsmutsade på grund av " Erikas " förlisning .
Var och en vet att ju mer tiden går desto större blir risken för att denna allvarliga olycka upprepas .
Den amerikanska lagstiftning , som antogs 1990 till följd av " Exxon Valdez " grundstötning på Alaskas kust , förbjuder tillträde till amerikanska hamnar för oljefartyg som inte uppfyller de stärkta och strängt kontrollerade säkerhetskriterierna .
Resultatet blir oundvikligen att de oljefartyg som inte uppfyller kriterierna kommer att dras - mer och mer - till europeiska vatten , vilket därmed ökar de troliga föroreningsriskerna .
Europaparlamentet måste således i första hand ta itu med dessa problem och först hos Europeiska kommissionen och därefter hos medlemsstaternas regeringar utan dröjsmål få till stånd att en mängd bestämmelser införs för att skydda havs- och turistverksamheterna vid den europeiska kusten .
Det är nödvändigt att utan dröjsmål inrätta en operativ europeisk maritim byrå vars främsta mål skulle vara att enligt normaliserade och enhetliga metoder samordna säkerhetskontroller på oljefartyg som anlöper europeiska hamnar .
Kära kolleger , att utarbeta och rösta fram en resolution är otvivelaktigt nödvändigt men det viktiga just nu är att vidta konkreta , kraftiga och modiga åtgärder som kan förhindra nya katastrofer .
Gemensam resolution om stormar i Europa .
( FR ) Den storm som har drabbat Europa och i synnerhet Frankrike påkallar för min del flera kommentarer och iakttagelser : 1 - Även om det inte är odiskutabelt fastställt att det finns en länk mellan denna storm , växthuseffekten och föroreningen är dessa händelser åtminstone en varning för vad som skall komma i framtiden om vi fortsätter att förorena vår planets atmosfär på ett oöverlagt sätt .
2 - Även om man i Europa också ofta har byggt billigt och föredragit elektriska luftledningar , som ofta är mycket fula visuellt mäter vi för närvarande de reella och tunga kostnaderna av dessa felaktiga besparingar .
3 - I de åtgärder som vidtagits för att reparera stormens förstörelse har vi kunnat konstatera både våra svagheter och vår brist på medel samt på samma gång de starka solidaritetskänslor som visats och den lika stora betydelsen av offentlig tjänst i vissa av våra offentliga företag som ofta har förtalats av den dominerande ultraliberala ideologin .
Jag vill hylla samtliga anställda och personalen i de företag som har arbetat ihärdigt och generöst för att återupprätta trafiken , återställa elektricitet och telefon samt hjälpa till med att skaffa nya bostäder åt de katastrofdrabbade familjerna .
4 - Om EU avslutningsvis vill förbli eller stå medborgarna nära måste man ingripa med betydande finansiella medel .
Dessutom måste medlemsstaterna , som ofta är överdrivet försiktiga , ge EU de nödvändiga finansiella medlen . .
( FR ) Problemet med stormarna , som olika europeiska länder har haft , visar hur ömtåligt vårt samhälle är , som likväl präglas av sin ekonomiska och tekniska utveckling .
Vi inser att vi inte är skyddade från de katastrofala konsekvenser som katastrofer av klimatologisk art , såsom översvämningar , jordbävningar eller jordskred , kan medföra .
Vissa länder har kunnat lösa problemet med ersättning åt offer för sådana fenomen .
Frankrike är ett exempel därpå , men det är ett stort land med betydande resurser .
Så är inte fallet för mindre länder .
I Belgien är således ett projekt för ersättning åt offer för naturkatastrofer i gång sedan tio år tillbaka .
Det är på europeisk nivå som de olika projekten har råkat i konflikt .
Först och främst , även om det var möjligt före genomförandet av den inre marknaden att föreskriva priser och självrisker , är det inte längre så och det verkar för mig vara normalt .
Däremot är det svårare att gå med på att det inte är möjligt att planera upprättandet av en ömsesidig kassa för återförsäkring , hos vilken de företag som är verksamma på den belgiska marknaden skulle tvingas försäkra sig .
Sedan skulle statens garanti bara kunna gälla om systemet har förbrukat samtliga medel ( med antagande av att en större katastrof inträffar ) .
Vi har dock en prioritering : att erbjuda katastrofdrabbade en total obegränsad garanti .
Ödet har redan kastat sig över dem utan att de är ansvariga , måste de få ytterligare svårigheter genom ett alltför svagt försäkringsskydd ?
Statens garanti är därför absolut nödvändig , eftersom ingen traditionell återförsäkring ger dem obegränsade villkor .
Det är enda sättet att ha ett lagom pris för konsumenten .
Begäran om en klassisk återförsäkring kommer att få en regleringseffekt på världsnivå , vilket betyder att de belgiska försäkringstagarna kommer att någonstans betala Centralamerikas orkaner ...
Tanken är inte att ta avstånd , utan att skaffa ett rättvist system , som är skyddat från att vara beroende av marknadslagarna .
Jag vill tillägga att det är enda sättet för staten att få garanti för att systemet fungerar med respekt för det allmänna intresset , samtidigt som man håller ett öga på anhopningen och användningen av tekniska bestämmelser .
Om denna insynsrätt inte tillåts kommer staten aldrig att gå med på att lämna garanti .
En kontrollerad återförsäkringsmekanism är det enda som gör det möjligt att undvika att riskerna väljs av marknadens naturlagar .
Om en nationell solidaritetsmekanism inte garanteras av ett system , som undantas till och med temporärt från marknadslagarna , kommer de dåliga riskerna att uteslutas medan det är just de riskerna som man försöker skydda ( t.ex. : bostäder vid flodstränder ) .
Därför ställer jag frågan om ett undantag från europeisk rätt , från den klassiska konkurrensrätten .
Det är för övrigt en tanke som är förenlig med fördraget .
I artikel 87.2 tillåts statliga stöd " för att avhjälpa skador som orsakats av naturkatastrofer " .
Sannolikheten för att sådana katastrofer upprepas är långt ifrån osannolik .
Lösningar bör också hittas för att finansiera skadeersättning åt offer för naturkatastrofer .
Ett temporärt undantag från konkurrensrätten skulle ge ett hopp om att lösa detta oroväckande problem i ett land som Belgien . .
( FR ) Jag röstade självfallet för resolutionerna om stormar och oljeutsläpp och jag vill framföra mitt deltagande till de drabbade befolkningarna .
Jag tänker särskilt och med värme på invånarna i min region , Champagne-Ardennes , som drabbades hårt av stormarna i december .
Jag beklagar de nya konsekvenser som oljeutsläppen skulle kunna få för kommunerna utmed Atlantkusten .
Jag oroar mig över vilka möjligheter som kommer att finnas kvar för båthamnar och lokala myndigheter att erövra den blå flaggan 2000 .
Den blå Europa-flaggan vittnar sedan 20 år om kommunernas avsevärda ansträngningar för att uppmuntra en ekonomisk utveckling som tar hänsyn till miljön .
Ett femtiotal kommuner i de 5 departement som drabbats av oljeutsläppen berörs av den blå flaggan 2000 .
Jag oroas också av rykten om en begäran att skjuta upp tilldelningen av blå flaggor till de franska stränderna vid Atlanten .
Vad skall man då säga om strändernas förlorade goda rykte , om orättvisan , eftersom vissa kommuner inte längre skulle ha någon flagga medan andra fortfarande har det .
Skall man acceptera att den ges till några kommuner för att förbättra en hel kusts rykte inför turisterna , eller inte ge den till någon av dem för att få viss rättvisa ?
Jag ber staterna och Europeiska unionen att lindra svårigheterna som uppstått på grund av dessa katastrofer , genom att lämna långfristigt ekonomiskt stöd , naturligtvis , men också genom ett " moraliskt " stöd ( - dessa resolutioner bidrar till detta - ) till de befolkningar som skadats in i själen av nedsmutsade stränder , uppryckta träd och skogar som jämnats med marken och förstörts .
Tidsbegreppet är viktigt för vi talar inte , som de multinationella företagen , om kortfristiga åtgärder , som de multinationella företagen , utan om århundraden för att återplantera Frankrikes skog , och det är en lektion i blygsamhet .
Gemensam resolution om fredsprocessen i Mellanöstern Herr talman !
Jag har i förväg anmält att jag vill avge en röstförklaring angående resolutionen om fredsprocessen i Mellanöstern .
Europaparlamentet har tidigare uttalat sitt stöd för en palestinsk stat och upprepar detta i punkterna 2 och 3 i dagens resolution .
Som svensk kristdemokrat anser jag att Europeiska unionen kan lämna ett bidrag till en bestående fred i Mellanöstern , ytterst baserad på demokrati , politisk pluralism , respekt för mänskliga rättigheter , rättsväsendets oberoende samt en social och ekologisk marknadsekonomi .
Detta kan ske genom att EU agerar på ett sådant sätt att det väcker mer förtroende och tilltro än i dag hos befolkningen i Israel , Mellanösterns enda demokrati .
Att därför i punkterna 2 och 3 nämna frågan om ett eventuellt bildande av en palestinsk stat bidrar inte till en sådan förtroendeskapande process .
Den amerikanska statsledningen har aldrig uttalat sig för en palestinsk stat , men äger samtidigt ett stort förtroende i regionen som fredsmäklare med konstruktiva bidrag .
En sådan roll skulle även Europeiska unionen kunna ikläda sig .
Dagens uttalande om en palestinsk stat stärker inte EU : s framtida möjligheter att göra detta .
Därför har jag i slutomröstningen lagt ned min röst . .
( IT ) De senaste nyheterna från Tel Aviv visar att fredens vägar , till skillnad från försynens , dessvärre inte är oändliga .
De kan blockeras och störas av terrorattacker , de kan fyllas av oskyldiga offer , de kan avbryta eller bromsa ansträngningarna från de människor av god vilja , på ena eller andra sidan , som uppriktigt önskar skapa fred .
Avtalet från Sharm el-Sheikh och förhandlingarna i Shepherdstown visar att , trots de skilda utgångspunkterna , så kan man komma fram till kompromisser på vägen mot det fredsmål som tyvärr fortfarande inte kan skönjas .
Det döljs av attentatens rökridåer , bojkottas av terrorister , fjärmas av fundamentalister av olika slag , personer som alltid är fiender till stabilitet och säkerhet .
För det är just säkerheten som är en av de grundläggande faktorerna när det gäller om vi skall lyckas : utan säkerhet kan det inte finnas någon fred , och utan fred i Mellanöstern kommer Medelhavet att förbli ett osäkert område , vidöppet för alla slags äventyrligheter .
Å andra sidan är den israeliske premiärministern Baraks inställning fullt begriplig , när han föreslår att den palestinska presidenten Arafat med en eller två månader skall skjuta upp den tidsfrist som satts till den 13 februari för att sluta ett ramavtal om de viktigaste punkterna i den framtida permanenta statusen för det palestinska territorium som Israel ockuperar sedan 1967 .
Även den uppskjutna tredje ronden i fredsförhandlingarna mellan Israel och Syrien omfattas av detta klimat av osäkerhet , en osäkerhet som beror på att det inte finns någon garanterad säkerhet .
Å andra sidan är vi övertygade om att fastställandet av en ny gräns mellan Israel och Syrien , en gräns som förutsätter en fredlig lösning av frågan om Golanhöjden och som tar hänsyn till båda ländernas behov av säkerhet , är ett nödvändigt villkor för att skapa nya fredliga relationer mellan de berörda folken och för att avlägsna riskerna för nya attentat och det våld som skulle bli följden .
Att sluta nya fredsavtal mellan Israel och Syrien ligger i hela Medelhavsområdets intresse och det skulle utgöra ett icke ringa bidrag till upprättandet av en ny balans i Mellanöstern .
Vi är alla övertygade om att det i världen även finns och opererar , ibland med en oerhörd grymhet , personer som motsätter sig balans och säkerhet .
Det är dessa personer som är fredens verkliga fiender .
De utnyttjar alla upptänkliga medel för att destabilisera regeringar och skapa oordning .
De finns i de områden där det råder spänningar , i själva verket provocerar de många gånger fram spänningar medvetet för att avbryta förhandlingar eller för att underblåsa stämningar bland allmänheten i syfte att utöva påtryckningar på regeringarna .
Europa måste ha modet att avslöja dessa krafter och att erbjuda sina tjänster , inte bara som medlare eller rådgivare på diplomatisk nivå , i fredsprocessen , utan även när det gäller att agera med auktoritet och kraft gentemot fredens fiender .
Det är otänkbart att de förbindelserna hela tiden skall ödeläggas av våld och attentat .
Terrorismen - för det är detta det handlar om - måste alltid fördömas och bekämpas .
Vi står nära våra israeliska vänner varje gång de drabbas av blind och avskyvärd terrorism , men vi måste också hela tiden bli effektivare i kampen mot dem som sätter vapen i händerna på terroristerna .
Om inte vägarna till fred kan bli oändliga , så måste vi se till att åtminstone de vägar är det som leder till att vi stoppar och oskadliggör dessa dödens handelsmän , dvs. de som är fredens verkliga fiender .
Resolutioner om skatt på kapitalrörelser Herr talman !
Europaparlamentets resolution om internationella kapitalrörelser som vi just förkastade , tog upp ett stort och intressant ämne men behandlade det tyvärr på ett ytligt och slarvigt sätt .
Uppriktigt sagt förtjänade ämnet bättre .
Efter några osammanhängande beaktanden avslöjade resolutionen i punkt 9 sitt verkliga syfte , nämligen att begära att " kommissionen inom sex månader skall upprätta en rapport rörande intresset och genomförbarheten av en skatt på internationella spekulativa kapitalrörelser " .
Om man tar upp frågan från den synvinkeln är jag ledsen att säga att det inte fanns någon grund för den begärda rapporten .
Alla vet redan att det är omöjligt .
Det är nämligen fullständigt omöjligt att skilja en spekulativ kapitalrörelse från en icke-spekulativ kapitalrörelse , om man inte använder godtyckliga och byråkratiska kriterier som skulle snedvrida handelsutbytet .
Och även om man lyckades med det , måste man ändå skilja de goda spekulationerna , som siktar till att ifrågasätta konstgjorda situationer för att i högre grad ta hänsyn till den reella ekonomin , från de dåliga spekulationerna , om vilka man skulle föreskriva , också godtyckligt för övrigt , att de huvudsakligen siktar till att skada andra .
Detta angreppssätt skulle vara ännu omöjligare än det föregående .
Kort sagt Europaparlamentets resolution var i denna form fullständigt utanför ämnet .
Problemet hade dock kunnat formuleras på ett annat sätt .
Man hade kunnat undra om det var lämpligt att införa en skatt på samtliga internationella kapitalrörelser , vilka de än är , utan att ge sig in på att göra omöjliga skillnader .
Det är en mer sansad fråga , men än en gång ställdes den inte .
På den andra frågan svarar jag likväl att en sådan enhetlig skatt troligen inte skulle lösa de valutakriser som oftast beror på verklig bakomliggande obalans .
I stället för att införa en ny skatt för att för övrigt mata kassor , om vilka vi inte vet någonting , skulle det var bättre att sanera den ekonomiska politiken och dra ner befintliga skatter och avgifter , i synnerhet på arbete . .
( EL ) Jag tycker att det är positivt att frågan om beskattning av de internationella kapitalrörelserna äntligen har kommit upp till diskussion och beslut i Europaparlamentet .
Det var ett välkommet initiativ från vår grupp , Europeiska enade vänstern , som sedan har fått stöd även av andra grupper .
Problemet är särskilt stort , om vi betänker att transaktionerna på aktiemarknaderna runt om i världen dagligen uppgår till 1 800 miljarder dollar och att den årliga handeln med varor och tjänster är i storleksordningen 6 000 miljarder dollar , vilket alltså motsvara fyra dagars spekulativ aktiehandel .
Ordförande Delors hade rätt , när han liknade den globala ekonomin med ett kasino .
Det är positivt att parlamenten i Finland och Kanada har uttalat sig för kapitalbeskattning , liksom även FN : s konferens för handel och utveckling ( UNCTAD ) i Förenta staterna .
Kommissionen måste lägga fram ett förslag om att införa en skatt på de kortfristiga kapitalrörelserna av spekulativ karaktär , av samma typ som Tobinskatten , liksom det portugisiska och det franska ordförandeskapet måste placera frågan bland sina prioriteringar .
En sådan skatt , låg men progressiv , måste vara utformad på ett sådant sätt att den inte får negativa följder för realekonomin - handel och investeringar - och så att den gör det möjligt att säkerställa medel till utbildningen , miljön eller tillväxten .
Denna åtgärd måste utgöra ett första steg mot att utforma ett regel- och skattesystem med vilket vi kan bemöta fenomenet med den internationella spekulationens enorma tillväxt .
Jag röstade för det gemensamma resolutionsförslaget , men det är beklagligt att att kristdemokraterna och liberalerna inte tillät att det röstades igenom . .
( DA ) Vi har röstat för kompromissförslaget mot bakgrund av de sunda avsikter som uttrycks .
Men samtidigt måste det påpekas att det är av avgörande betydelse att diskussionen om införande av en eventuell Tobinskatt sker på en global nivå vid internationella och nationella fora , och utan att det som bieffekt ökar EU : s behörighet på bekostnad av dessa . - ( FR ) Vårt ekonomiska system har visat sina gränser .
Finanssfären är inte i fas med den reella ekonomin och rubbar den alltför ofta .
Den höga arbetslösheten i våra länder , ökningen av klyftan mellan norr och söder samt den ökade fattigdomen i hela världen vittnar om den tråkiga verkligheten .
Världsomfattande kapitalrörelser är destabiliserande !
Därför måste vi söka efter åtgärder i syfte att beskatta transaktionerna på valutamarknaden så att vi gör dem mindre flyktiga och förhindrar kortsiktiga spekulativa operationer .
En skatt såsom den som James Tobin , Nobelpristagare i ekonomi , tänkt ut skulle utgöra ett sandkorn i spekulationens alltför väloljade kuggar och de stora summor som den skulle kunna frigöra är goda argument för att den skall tillämpas , när man vet att även om man sätter en mycket låg sats ( omkring 0,05 procent ) skulle den inbringa nära sexhundra miljarder franc varje år enligt de mest pessimistiska uppskattningarna !
Förenta nationernas konferens om handel och utveckling ( UNCTAD ) föreslår därför att denna summa skall återbetalas till de stater , i vilka skatten skulle tas ut , samt till en omfördelningsfond för de fattigaste länderna .
Denna rikedom som således skulle tas ut från de stora internationella kapitalisterna skulle omfördelas till medborgarna och skulle kunna utgöra en enorm drivkraft för utveckling i de minst gynnade länderna .
Vi skulle äntligen befinna oss i en logisk situation där solidariteten skulle ersätta egoismen .
Av samtliga dessa skäl röstade jag för resolutionen och jag är glad att kammaren återupptagit ärendet med risk för att stöta sig med samvetslösa spekulatörer som genom sina handlingar destabiliserar de känsligaste ekonomierna och ibland till och med vårt system i sin helhet , såsom finanskriserna i Sydostasien nyligen vittnar om . .
( FR ) Vi har röstat för begäran om att debatten om Tobinskatten skall sättas upp på föredragningslistan eftersom vi är övertygade om att dess , till och med begränsade , tillämpning i Europa skulle vara ett första steg till större social rättvisa och en annan fördelning av rikedomar .
Vi gör oss ändå inte den minsta illusion om att denna skatt ensam skall kunna avskaffa själva orsakerna till den fattigdom som är förbunden med det ekonomiska och finansiella system som dominerar världen .
Vi röstar för allt som siktar till att uppmana kommissionen att granska Tobinskattens genomförbarhet .
Vi röstar däremot inte för ingresserna i kompromissresolutionen från socialdemokraterna , den europeiska enhetliga vänstern , de gröna och de liberala , som siktar till att försvara och reglera det dominerande ekonomiska systemet och " säkra de globaliserade finansmarknadernas funktion , till och med om de blivit befriade från sina överdrifter " . .
( FR ) De valda från arbetarkampen kommer att rösta emot kompromissresolutionen om beskattning av kapitalrörelser .
Under en både futtig och utopisk förevändning av att " stabilisera " det internationella finansiella systemet och " befria det från sina överdrifter " påpekas det framför allt i resolutionen att målet är att bevara det .
Vår synvinkel är att mänskligheten inte bara skall befrias från överdrifter i det finansiella systemet i världen utan från det finansiella systemet själv och från den kapitalistiska organisationen av ekonomin , varav det är en väsentlig beståndsdel .
Det är inte bara det kortsiktiga spekulativa kapitalet på finansmarknaderna som utgör ett ofantligt , materiellt , socialt och mänskligt slöseri för samhället utan kapitalet rätt och slätt .
De permitteringar och indragningar av arbetstillfällen som pågår , från Michelin till Alsthom , som nästan samtliga storföretag , som likväl är lönsamma , i Europa genomför endast i syfte att få aktiekursen att stiga på börsen : är det spekulation eller kapitalets normala verksamhet ?
Om en resolution tydligt föreslog att Tobinskatten skulle införas , hade vi inte röstat emot för att vår röst inte skall blandas samman med rösterna från det kapitalistiska systemets självbelåtna beundrare som ser skatt på storkapitalet såsom en förolämpning .
För vår del är det politiska mål som vi föreslår arbetarklassen att den inte bara föreskriver mycket stora skatter på det spekulativa kapitalet , utan också på alla kapitalistiska storföretags vinster samt på den rika klassens privata förmögenheter så att de pengar som således kommer att koncentreras i statens händer skall kunna tjäna till att skapa nyttiga arbetstillfällen i offentlig tjänst .
Men den löjligt låga Tobinskatten är visserligen inte ett mått på social rättvisa , den skulle inte ens störa spekulanterna , och i stället för att sätta upp hinder för den kapitalistiska ekonomins slöseri och orättvisa skulle den bara tjäna till att dölja det . - ( PT ) Den oro som visas i förslaget till gemensam resolution är mycket viktig , och tar upp ett allvarligt problem och vi får inte fortsätta att stoppa huvudet i sanden inför det och låtsas som om det inte existerar .
Jag stödde därför uttryckligen samtliga punkter i det gemensamma resolutionsförslaget , utom punkterna 4 och 8 , där jag avstod därför att de gick in på speciella egenskaper som var onödiga eller ofärdiga .
Punkt 4 därför att jag inte tycker att en lätt analys av ett mycket komplext problem är korrekt i någon betydelse av ordet , punkt 8 därför att det rekommenderade omedelbara åtgärder mot off-shore-centren , vilket avskilt från en allmän och balanserad ram skapar en ömtålig situation i Portugal vad gäller nuvarande off-shore på Madeira .
Eftersom denna punkt 8 emellertid antogs av en majoritet - såg jag mig tvungen , mot min vilja , att avstå även i den allmänna slutomröstningen .
Jag beklagar att den gemensamma resolutionen inte antogs , då det är bråttom att ta upp denna fråga i mer försiktiga ordalag , men med rätt inriktning .
Jag stödde därefter inget resolutionsförslag från de olika grupperna , vilka vi röstade om var för sig , eftersom inget av dem innehöll den balans som det gemensamma resolutionsförslaget försökte uppnå .
Betänkande ( A5-0096 / 1999 ) av Cunha Herr talman !
Även när det gäller detta betänkande som avser en utvärdering av fiskeriprogrammen , är jag som företrädare för Pensionärspartiet positiv .
Det måste vara riktigt att ha sanktioner för dem som inte tillämpar direktiven , men jag måste också säga att min röstförklaring i kammaren fredagen den 17 december 1999 , dvs. under förra seklet , nådde ända fram till fiskarna själva , som - eftersom de , som vi alla vet , inte kan tala - skriftligen meddelat mig följande : " Bra , du talade i vår sak !
Tala nu också för oss småfiskar , framför allt eftersom du själv är en liten fisk , men tala också för de gamla fiskarna , de som skulle vilja leva länge och som därför ser positivt på att man begränsar fisket på de platser där det råder brist . "
De ber mig också - men det skall jag göra i ett annat sammanhang - att lägga fram deras förslag när det gäller måtten på fiskenäten så att de skall kunna leva länge och även de en dag bli pensionerade fiskar . - ( PT ) Min röstning sammanfaller med Portugals folkparti CDS - Partido Populars ståndpunkt i denna fråga : å ena sidan är vi starkt kritiska mot den gemensamma fiskeripolitiken , vilken har lett till så stora skador för fisket och fiskarna i Portugal , och vi ser med särskild misstänksamhet på kommissionär Fischlers agerande , å andra sidan stöder vi ståndpunkterna i Cunhas betänkande och kräver effektiva kontroll- och övervakningsåtgärder från kommissionens sida - kommissionen diskriminerar tilläggsvis de länder som , såsom Portugal , uppfyller målen då man inte verkligen straffar de länder som inte uppfyller dem .
Jag röstade således för de första och sista delarna i punkt 6 , även om jag lade ner min röst angående dess mellanpassager som rekommenderar en konkret sanktion - , dels för att det är för tidigt innan det finns en lämplig rättslig grund , dels för att en sådan ekonomisk sanktion skulle kunna vara olämplig i andra situationer , när det bara handlar om brott mot föreskrifter .
Jag lade också ned min röst i den allmänna omröstningen , dels för att just dessa sista passager antogs , dels för att punkt 5 inte blev föremål för en separat omröstning .
Även om CDS-PP stöder den oro som visas i betänkandet och resolutionen vill det inte för närvarande stödja något som kan tolkas som ett stöd för en gemensam fiskeripolitik som i praktiken har lett till skadliga effekter för Portugal .
Herr talman !
En ordningsfråga .
Jag vill tala om hur glad jag är att se er på er plats i en sådan god form efter er sjukdom nyligen !
Tack så mycket !
Jag förklarar omröstningen avslutad .
( Sammanträdet avbröts kl .
12.44 och återupptogs kl .
15.00 . )
 
DEBATT OM AKTUELLA OCH BRÅDSKANDE FRÅGOR Nästa punkt på föredragningslistan är den aktuella och brådskande debatten om frågor av större vikt .
 
Tjetjenien Vi börjar med den gemensamma debatten om följande resolutionsförslag om Tjetjenien : ( B5-0048 / 2000 ) av Schori och Krehl för PSE-gruppen om situationen i Tjetjenien , ( B5-0065 / 2000 ) av Haarder m.fl. för ELDR-gruppen om Tjetjenien , ( B5-0067 / 2000 ) av Markov m.fl. för GUE / NGL-gruppen om kriget i Tjetjenien , ( B5-0080 / 2000 ) av Schroedter m.fl. för Verts / ALE-gruppen om kriget i Tjetjenien , ( B5-0082 / 2000 ) av Oostlander m.fl. för PPE-DE-gruppen om situationen i Tjetjenien .
Herr talman , mina damer och herrar !
Ännu en gång är det med rätta som parlamentet befattar sig med läget i Tjetjenien .
Under tidigare sammanträden har vi gång på gång betonat vikten av att den ryska federationen finner en fredlig och politisk lösning på problemet .
Vi har verkligen vädjat till den ryska regeringen om att inte agera på ett sätt som skadar samtliga internationella konventioner som man har skrivit under .
Tyvärr kan vi ännu inte rapportera om någon avspänning i kriget .
Mycket värre än så !
Situationen har förvärrats avsevärt .
Situationen för civilbefolkningen i Tjetjenien har blivit outhärdlig .
Vi har ingen möjlighet att vidta humanitära åtgärder , trots att vi vid upprepade tillfällen har understrukit och den ryska federationen åtminstone på toppmötet i Istanbul har försäkrat att det skall bli möjligt för såväl observatörer från OSSE som för humanitära organisationer att komma till Tjetjenien .
Jag har inget annat val än att upprepa det som redan har sagts här i kammaren och som vi ännu en gång vill understryka i ett gemensamt resolutionsförslag .
Vi vill få till stånd en politisk lösning på konflikten .
Här måste alla parter uppmanas att delta i förhandlingar .
Vi vill underlätta situationen för civilbefolkningen genom att återigen uppmana den ryska federationen att acceptera att humanitära organisationer bereds tillträde till Tjetjenien och även att släppa in observatörer från OSSE i Tjetjenien .
Herr talman !
Kriget i Tjetjenien började till stor del på grund av skäl som mer har att göra med den ryska inrikespolitiken än med situationen i själva Tjetjenien .
Jag fruktar därför också att det inte finns mycket hopp om att kriget skall sluta förrän Putin vunnit valet den 26 mars eller möjligen tidigare genom en total rysk seger i kriget .
Det viktiga är vad som händer när konflikten äntligen är förbi och det är svårt att förutse .
Det är tydligt att problemen i Tjetjenien och i norra Kaukasus , som hör till de fattigaste områdena i Ryssland , inte är över när själva kriget tar slut .
När den tjetjenska befolkningen kan återvända till sitt land kommer de att återfinna mycket litet som de kan bygga upp sin existens med igen .
Efter det förra kriget blev det ingenting av den utlovade ryska återuppbyggnaden och det var svårt att erbjuda utländsk hjälp på grund av problem både från rysk och från tjetjensk sida .
Samtidigt är det också bra att titta på positiva exempel , till exempel de framsteg som gjorts i de tre oberoende kaukasiska staterna , Armenien , Azerbajdzjan och Georgien .
Där finns det inget krigshot längre och de europeiska institutionerna måste känna till hur situationen är där .
Så kan det nämligen också se ut .
Herr talman !
Kriget i Tjetjenien har nu rasat i fyra månader .
Europaparlamentet har fördömt det , krävt vapenstillestånd samt att den politiska dialogen skall öppnas .
Parlamentet har bidragit till att humanitär hjälp ges och att ekonomiskt stöd från Europeiska unionen också styrs om i den riktningen .
Något slut på kriget och på civilbefolkningens lidanden är inte inom synhåll , än mindre en hållbar lösning på konflikten .
Har EU verkligen gjort allt som står i dess makt ?
Faktum är att rådet och vissa medlemsländer , däribland även Tyskland , är utomordentligt återhållsamma vad beträffar politiska , diplomatiska och ekonomiska reaktioner på Rysslands oavlåtliga vägran att delta i den politiska dialogen .
Europeiska unionen och dess medlemsländer måste tydligt visa att denna fullkomligt överdrivna användning av militärt våld för att lösa konflikten i Tjetjenien och den massiva kränkningen av mänskliga rättigheter inte är acceptabla .
Europaparlamentet bör kämpa för att få partnerskaps- och samarbetsavtalet med Ryssland upphävt tills Ryssland accepterar ett vapenstillestånd .
Dessutom bör vi uppmana medlemsländerna att vidta kompletterande politiska , diplomatiska och ekonomiska sanktionsåtgärder .
Vapenaffärer liksom det finansiella stödet till de krigförande parterna måste omedelbart stoppas .
Rysslands suveräna rätt att skydda sin territoriella integritet och att förfölja terrorism är obestridlig .
Frågan är med vilka instrument man gör detta .
Förhållandet mellan dialog och samarbete med Ryssland och sanktioner med hänsyn till kriget är en komplicerad balansgång .
Vi får inte förödmjuka och isolera Ryssland , vilket har varit fallet många , många gånger under de gångna decennierna .
Det ömsesidigt fördelaktiga samarbetet och partnerskapet med Ryssland är oundgängligt för en fredlig utveckling i Europa .
Europeiska unionens utrikespolitik är dock trovärdig endast om man i samband med krig och massiva kränkningar av de mänskliga rättigheterna inte drar sig för att vidta konsekventa politiska , diplomatiska och ekonomiska åtgärder .
Herr talman !
I går menade mina kolleger att Tjetjenien har stått som nummer 1 på föredragningslistan om och om igen i flera månader nu .
Och vad har kommit ut av alla våra krav ?
Vi måste - som Sakellariou ju mycket tydligt sade - hela tiden upprepa våra krav .
Inte heller jag anser att vi får tröttna , för så länge det militära våldet mot den egna civilbefolkningen i Ryssland verkligen ökar dramatiskt måste vi höja våra röster och säga : " Nu är det nog !
Detta accepterar vi inte !
Detta är en kränkning av internationella mänskliga rättigheter !
Detta är ingen intern angelägenhet för Ryssland . "
Listan över krigsförbrytelserna blir allt längre .
Det må gälla ungdomarna som tillfångatogs i flyktingkolonnerna , det må gälla listan över de många våldtäkterna , vilken anlände till mitt kontor i dag och som har sammanställts av oberoende observatörer för de mänskliga rättigheterna .
Kvinnorna i det islamiska samhället försätts ju härigenom i en mycket dramatisk situation .
Därför måste vi ta oss an dem alldeles särskilt .
Det är just de många små enskilda ödena som uppmanar oss att inte tiga .
Många viktiga dricksvattenreservoarer har på grund av bombningarna börjat förgiftas av olja .
Jag ber mina kolleger att godkänna detta ändringsförslag .
Det nådde oss efter det att vi gemensamt hade diskuterat resolutionen .
Vi kan helt enkelt inte bara sitta och titta på !
I motsats till Kosovo är det faktiskt så att de 100 000 flyktingarna är utan internationell hjälp i Ingusjien .
Denna pyttelilla grannrepublik är totalt överlastad .
Jag måste säga att jag egentligen är förvånad över att vi över huvud taget inte får något svar på våra krav från kommissionen .
Jag väntar mig i dag egentligen en något mer konkret beskrivning av hur ni följer parlamentsbesluten och besluten från Helsingforsresolutionen .
Vad ni hade att komma med i går var verkligen en skam gentemot parlamentet !
Vidare förväntar jag mig en undersökning av huruvida det som sker i Ryssland verkligen är förenligt med artikel 2 i ...
( Talmannen avbröt talaren . )
Herr talman !
Den ryska federationens regering ser sig själv som en fullvärdig medlem av till exempel Europarådet .
Det medför skyldigheter som sträcker sig mycket längre än till diverse internationella avtal för skydd av de mänskliga rättigheterna , mycket längre än krigsrätten .
De förbindelser som vi ingått med Ryssland i olika fördrag pekar också i den riktningen .
Det sätt som den ryska regeringen försöker lösa sina problem med Tjetjenien på strider dock helt och hållet mot de internationella reglerna .
Vi kan föreställa oss att man var tvungen att reagera mot till exempel terrorism och aggressioner gentemot Dagestan .
Det är så att myndigheterna i Tjetjenien inte hur som helst kan ses som företrädare för en reglerad demokratisk rättsstat .
De kunde till exempel inte förhindra de brutala kidnappningarna och gisslandramerna på det egna området .
De medel som Ryssland använder är dock oproportionella och bör fördömas i sig , och därvid menar jag särskilt bombningarna av befolkningen och behandlingen av den del av befolkningen som håller på att lämna landet .
Vi är skyldiga att motsätta oss det .
Inte av självgodhet , eftersom jag själv kommer från en före detta kolonialmakt så känner jag nämligen till den sortens krig och den ånger över begångna missdåd som kommer upp till ytan först tjugo , trettio år senare .
Framtiden för Ryssland och Tjetjenien rör oss dock i hjärtat och därav denna uppmaning .
Vi stöder därför också den här resolutionen av hjärtat .
Resolutionen riktar främst in sig på humanitära aspekter , på ekonomiska bidrag , på en förflyttning av Tacis-programmet i den riktningen , på diplomatiska förhandlingar och möjligtvis på förhandlingar inom ramen för OSSE angående stabiliteten i Kaukasus .
Vi i Europeiska unionen vill samarbeta med internationella organisationer som Ryssland vill ha och förväntar sig stöd ifrån .
I varje fall måste vi även på det här sättet , även med hårdhet om det är tvunget , fortsätta dialogen med Ryssland på alla möjliga sätt .
Herr talman !
Vad är det som har förändrats under de fyra månader som vi har arbetat med denna fråga ?
För det första har Putins mjuka kupp ägt rum - mycket smidigt på nyårsaftonen vid millennieskiftet - vilken har gett honom en mycket mäktig position men också gjort honom till en av vår tids största politiska krigsprofitörer .
Jag anser likväl att han bör utnyttja den makt han nu har till att göra slut på vad general de Gaulle har kallat paix des braves , de tappras fred .
Det är nu så att han har chansen att få ett slut på detta mordiska krig , och det utifrån en position som är rätt stark .
Om han inte lyckas är det möjligt att han kommer att få se sina presidentdrömmar gå under i ett blodbad .
En andra väsentlig punkt : ytterligare något har förändrats , och det är situationen i den ryska offentligheten .
Tack och lov förekommer det kritik .
Det kommer kritik från soldatmödrarna , det kommer kritik från media , från människorättskämpar .
De är fortfarande i minoritet , men det visar att nu som då även det ryska folket har ett levande samvete och att vi inte får göra det ryska folket ansvarigt för ledningen .
Den tredje punkten : jag anser att man i Tjetjenien har visat en beundransvärd motståndsvilja , varför jag har stora problem med punkt fyra i vårt beslut , för jag förstår till fullo att man försöker skydda människorna i Tjetjenien från att bli offer i ett folkmord .
Jag menar att vi i Europeiska unionens namn äntligen måste utöva ett massivt politiskt tryck genom att ta itu med artikel 2 i partnerskapsavtalet , genom att även kommissionen och rådet äntligen börjar utöva konkreta påtryckningar , vilket parlamentet ända från början har gjort inom ramen för sina blygsamma möjligheter .
Vi måste som EU tala med en röst och får inte överlåta åt Europaparlamentet att tala i klartext .
Vad den humanitära hjälpen anbelangar är jag av den åsikten att vissa oberoende organisationer som redan har lyckats med konkreta hjälpinsatser får oss att skämmas .
Jag känner till en barnmatstransport som man nu har lyckats genomföra .
Men sorgligt nog lyckas inte kommissionen bygga upp motsvarande kanaler i de omgivande trakterna , och jag skulle verkligen vilja veta varför kommissionen inte lyckas med det .
Här måste det till konkreta humanitära hjälpinsatser mot folkmordet , för det som sker i Tjetjenien är ingenting annat än ett folkmord .
Herr talman , kära kolleger !
Det är inte bara under de senaste fyra månaderna i och med denna andra militära konflikt som vi här i kammaren har diskuterat problemet mellan de kaukasiska folken och Ryssland .
Det har vi mycket ofta gjort även tidigare .
Hittills har vi dock inte rönt någon framgång i den aktuella militära konflikten som gäller Ryssland mot det tjetjenska folket .
Det råder fortfarande inte fred i området , och trots att Europaparlamentet hela tiden har visat en mycket tydlig politisk ståndpunkt har vi ännu inte lyckats .
Jag tror att nya politiska möjligheter har öppnat sig för oss i Ryssland efter valen till duman och president Jeltsins avgång .
Jag anser att Europaparlamentet också måste försöka att , vid sidan av överläggningarna om vilka sanktioner som är meningsfulla , föra en politisk dialog med de ryska politikerna .
Duman är sammansatt på ett sätt som den aldrig tidigare har varit , och detta ger oss även en chans att finna politiska bundsförvanter för att få ett politiskt slut på den militära konflikten i Tjetjenien så att freden äntligen kan göra sitt intåg där .
Vi alla vet att de kaukasiska folkens problem inte på långt när är lösta ens när den militära konflikten väl är över .
Därefter behöver vi en politisk dialog .
Vi behöver ett politiskt samarbete , för konflikten har ju inte uppstått först i dag .
Den har uppkommit ur de kaukasiska folkens historia i och mot Ryssland och mot deportation och mot rysk ockupation .
Jag anser att det vore helt i linje med Europaparlamentets strävan om vi kunde finna allierade för en politisk dialog även när den militära konflikten är slut .
( Applåder ) Herr talman !
Vi är naturligtvis upprörda över det barbariska ryska ingripandet i Tjetjenien , och upprörda över att se hur Boris Jeltsin och hans gelikar har kunnat utnyttja dessa massaker för att det elände som deras politik har försatt det ryska folket i skall glömmas bort .
Morden i Tjetjenien ger nu röster i Moskva .
Men upprördheten kan inte bara sammanfattas med detta .
Hur skall vi tolka den medbrottsliga passiviteten från västmakternas sida , som vill vara förkämpar för humanitär och militär nödhjälp och som inte tvekat att bomba Irak och f.d.
Jugoslavien ?
Dessa makter kastar för närvarande ljuva blickar på den alkoholmaffia som styr Ryssland .
Vi kan påminna oss de entusiastiska talen av amerikanska och europeiska ledare som prisade Boris Jeltsin förtjänster .
Genom att solidarisera sig med den ryska regeringen har de gett förtur åt återupprättandet av marknadslagarna till nackdel för skydd av folkens rättigheter .
Vi måste upphöra med detta skamliga hyckleri och kräva ett omedelbart tillbakadragande av de ryska trupperna och rätt till självbestämmande , det vill säga det tjetjenska folkets oberoende .
Herr talman , herr kommissionär , kära kolleger , jag skulle här vilja hylla Dimitri Neverovsky , medlem av det transnationella radikala partiet , medlem av mitt parti , som har dömts till två års fängelse för vapenvägran och för att ha motsatt sig kriget i Tjetjenien .
Jag skulle också vilja hylla det transnationella partiets förkämpar som ensamma i Moskva har demonstrerat mot kriget i Tjetjenien .
Jag tror tyvärr att vi inte kan hylla , av de orsaker som Schroedter påminde om , vår kommissionsledamot , Poul Nielson , som på fyra månader inte har haft ett ögonblick för att bege sig till Tjetjenien och till området för att se till att Europeiska unionen åtminstone på det humanitära planet - jag talar här inte om det politiska planet - åtminstone på det humanitära planet bemöter den pågående tragedin på ett tillfredsställande sätt .
Jag tror att det är mycket allvarligt .
Jag hoppas att vi inom de närmaste dagarna till slut kommer att kunna se Nielson i Tjetjenien , i området , i Ingusjien och äntligen ta hand om flyktingarna .
Herr talman !
Två röster från tjetjenska kvinnor , flyktingar .
Första citatet : " Min son är 13 .
Om vi vänder tillbaka är jag rädd att ryssarna arresterar honom omedelbart och låter honom försvinna " .
Andra citatet : " Rysarna är inga befriare utan ockupanter .
Förut var det islamiterna som terroriserade oss .
I dag är det de ryska soldaterna som gör det . "
Slutet på blodsutgjutelsen i norra Kaukasus verkar inte alls vara i sikte .
Utan någon som helst tvekan säger den ryska premiärministern och tillförordnade presidenten , Vladimir Putin , till en officiell delegation från Europarådet att de inte skall grunda sin kritik mot Kremlins krig på propagandamaterial .
Nej , Moskva har mycket riktigt redan från början lagt ner mycket energi på att redigera publiciteten kring detta det andra tjetjenska kriget på några få år .
Det hjälper dock inte .
Berättelserna från den enorma skaran av tjetjenska flyktingar talar sitt tydliga språk .
Inte heller låter alla ryska politiker sig toppridas och skrämmas av Putin och dennes sufflörer .
Den reformvänliga presidentkandidaten Grigorij Javlinskij till exempel , säger utan omsvep att det är brottsligt att utnyttja ett krig för valändamål .
Javlinskij yrkar för en dialog med de Tjetjeniens ledare och befolkning .
Denna ryska besinningsfullhet förtjänar vårt stöd .
Det reella hotande alternativet är annars ett i det närmaste utsiktslöst gerillakrig .
Den här , politiskt balanserade resolutionen från Europaparlamentet försöker i varje fall förhindra detta skrämmande och farliga scenario .
Effekterna av den kan vi hur som helst mäta när Putins utrikesminister , Ivanov , besöker Europarådet i Strasbourg .
Herr talman , bästa kolleger !
Vi har pressat Ryssland till en politisk lösning i Tjetjenien .
Våra hot om sanktioner har inte lett till några resultat .
För att kunna påverka den politiska lösningen i Tjetjenien måste man enligt min mening inleda en politisk dialog med den ryska ledningen om detta , alltså med politiska medel för en politisk lösning tillsammans med den nya ledningen .
70 procent av dumans ledamöter är nya , och Ryssland har en ny tillförordnad president .
Denna tillförordnade president har uttryckt sin vilja till politisk dialog .
Han har redan träffat en delegation från Europarådet och samtalat med den under tre timmar .
Mitt förslag är att parlamentets delegation till Moskva explicit för att föra politiska samtal med den nya ledningen .
För det andra föreslår jag att kommissionär Christopher Patten , som ansvarar för yttre förbindelser , också skall inleda politiska samtal om läget i Tjetjenien .
Med politiska medel kan man påverka det politiska krig som det nu handlar om . .
( FR ) Herr talman , kommissionen stöder fullt och fast ett långsiktigt partnerskap med Ryssland , grundat på partnerskaps- och samarbetsavtalet och på den gemensamma strategin , i syfte att stärka säkerhet och stabilitet i Europa och inom en bredare ram .
I enlighet med parlamentets tydliga och klara ståndpunkt anser kommissionen att det skulle vara ett misstag att avbryta samtliga kommunikationskanaler .
Vi bör i synnerhet var i stånd att diskutera med ryssarna om vår djupa oenighet och vår stora oro inför situationen i Tjetjenien .
Europeiska rådet som samlades i Helsingfors sände ett mycket tydligt budskap om den kritiska situation som civilbefolkningen befinner sig i och att Ryssland bör följa humanitära rättsregler , i synnerhet i samband med det ultimatum som gavs åt Groznyjs invånare , det överdrivna utnyttjandet av våld och tvång utan åtskillnad mot civilbefolkningen , hindren för en säker och snabb transport av humanitär hjälp av hjälporganisationer samt bristen på verklig politisk dialog med de legitima tjetjenska myndigheterna .
Efter toppmötet i Helsingfors har situationen inte förbättrats .
Trots att ultimatum till Groznyjs befolkning inte verkställdes är vi mycket bekymrade för civilbefolkningens nödläge och i synnerhet för de personer som befinner sig i Groznyj som i en fälla .
Villkoren för att genomföra de humanitära åtgärderna är fortsatt svåra .
Ingen utväg syns ännu när det gäller den militära konflikten , eftersom de ryska styrkorna möter ganska starkt motstånd .
Interimspresidenten , Putin , talar hädanefter om en förlängd åtgärd .
Fruktan ökar för att grannen Georgien skall dras med av den ostadiga situationen .
Ordförandeskapet och kommissionen arbetar aktivt med att tillämpa slutsatserna från Europeiska rådet i Helsingfors , det vill säga att ompröva genomförandet av den gemensamma strategin , upphäva vissa bestämmelser i samarbetsavtalet och strängt tillämpa handelsbestämmelserna , planera att överföra Tacis-medel till humanitär hjälp samt dra ner Tacis 2000 till ett grundprogram med begränsad omfattning .
Dessa frågor kommer att diskuteras nästa måndag av utrikesministrarna vid sammanträdet av rådet för " Övriga frågor " .
Det är tydligt att vi inte nu kan föregripa resultatet .
Men jag kommer att se till att min kollega Chris Patten informeras om de frågor som tagits upp vid denna debatt så att han kan föra dem vidare till rådet .
Jag skulle slutligen vilja betona att förklaringen från Helsingfors har tagit sig uttryck i konkreta åtgärder , i vilka parlamentets synpunkter särskilt beaktas , det vill säga uppskjutandet av undertecknandet av det vetenskapliga och tekniska avtalet och den stränga tillämpningen av handelsbestämmelserna , till att börja med en åtgärd inom stålsektorn mot exportavgifter på icke järnhaltigt metallskrot .
Kommissionen har dessutom beslutat att inte be budgetmyndigheten på nytt överföra de anslag från programmet för livsmedelshjälp till Ryssland som inte användes förra året .
Herr talman , har kommissionär Nielson avgått ?
Vi hör aldrig talas om honom .
Patten , om det som berör honom , ja , men Nielson , ansvarig kommissionär för humanitära frågor är fullständigt frånvarande .
Vi skall inte debattera detta , men jag vet att det finns förmildrande omständigheter till varför Nielson inte kan vara här denna vecka .
Talmannen meddelade det från ordförandeskapet i måndags .
Hon sade att Nielson personligen hade skrivit till henne för att förklara varför han inte kunde vara i plenum denna vecka .
Herr talman !
Det hör ju till ordningen att man tillåts ställa en kort fråga till kommissionären .
Jag undrar bara konkret - eftersom frågan inte har besvarats - ges det humanitär hjälp , ja eller nej ?
Har hjälp alltså getts hittills , jag menar inte i framtiden , utan nu , konkret .
Jag kommer att tillåta kommissionären att svara om han vill , men det är inte normalt att ställa följdfrågor under den aktuella och brådskande debatten .
Det rör sig om debatter med snäva tidsramar .
Men om kommissionären vill ta ordet , är han välkommen att göra det . .
( FR ) Herr talman , Nielson har redan betonat svårigheterna med att transportera den humanitära hjälpen .
Problemet finns framför allt i det avseendet .
Jag förklarar den gemensamma debatten avslutad .
Omröstningen kommer att äga rum kl .
17.30 .
 
Elfenbenskusten Nästa punkt på föredragningslistan är gemensam debatt om följande resolutionsförslag om Elfenbenskusten : ( B5-0049 / 2000 ) av Carlotti och Sauquillo Pérez del Arco för PSE-gruppen om situationen i Elfenbenskusten , ( B5-0063 / 2000 ) av Van den Bos för ELDR-gruppen om Elfenbenskusten , ( B5-0068 / 2000 ) av Sjöstedt och Alavanos för GUE / NGL-gruppen om situationen i Elfenbenskusten , ( B5-0077 / 2000 ) av Rod m.fl. för Verts / ALE-gruppen om Elfenbenskusten , ( B5-0087 / 2000 ) av Novelli m.fl. för PPE-DE-gruppen om statskuppen i Elfenbenskusten .
Dåliga regeringar måste försvinna genom valurnan och inte genom en gevärspipa .
Det gäller också för Elfenbenskusten .
Det stora och berättigade missnöjet med den korrumperade Bedié-regimen rättfärdigar inte en statskupp .
Det handlar nu om att de nya makthavarna håller sitt ord och snabbt återställer demokratin , fastställer en grundlag och genomför fria val under internationell tillsyn senast i juni .
Det är också av stor betydelse att man gör något åt korruptionen .
Om den nya regimen inte håller sina löften så måste samarbetsavtalet med Europa upphävas .
Den nationella enhetsregeringen har mycket litet tid på sig för att återställa det internationella förtroendet .
Ju fortare den själv försvinner via valurnan , desto bättre .
Kompromissresolutionen om situationen i Elfenbenskusten kräver att den demokratiska legitimiteten återställs .
Men vad handlar det om ?
Från den otrevliga franska kolonialdominansen genom Houphouët-Boignys diktatur och den lika auktoritära som korrumperade regimen under Konan Bédié , fram till Gueis militärregim har befolkningen i Elfenbenskusten aldrig haft verkligt fria val eller demokratiska fri- och rättigheter .
Bakom de hycklande fraserna om demokrati , ägnar man sig i resolutionen framför allt åt återupprättandet av statsmyndigheten och säkerheten för tillgångar .
Vår solidaritet går till den förkrossande majoriteten av befolkningen i Elfenbenskusten , arbetare , arbetslösa och småbrukare som inte har några tillgångar och redan helt enkelt bara svårt att överleva .
De har alltid tvingats stå ut med statens repressiva myndighet , förutom diktatur och elände .
Jag vill också påminna om den franska statens ansvar , alla regeringar sammantagna , som inte bara har stött enpartiregimen i Elfenbenskusten utan har fört fram den såsom ett exempel på stabilitet eller rent av demokrati för Afrika i sin helhet .
Allt detta för att bevara de stora franska industrikoncernernas intressen , koncerner vars rikedomar växer där samtidigt som de utarmar landet .
Låt oss då sopa framför egen dörr , för om Gueis rena militärregim och Bédiés falska demokrati bör fördömas , bör stormakterna och deras stöd åt de fattiga ländernas diktaturer fördömas ännu mer .
( Applåder ) Herr talman , herr kommissionär !
För några månader sedan hörde jag här Johan Van Hecke i förfärande och berättigade ordalag fördöma den dåvarande regeringen som nu avsatts genom en statskupp .
Jag håller med de kolleger som säger att det inte är det rätta sättet .
I ett sådant land finns det väl ändå inte så många bra sätt att göra något sådant på .
Den här regimen var en dålig regim .
Nu hoppas vi att en process kan komma i gång , demokrati tycker vi nämligen inte bara är fria val .
Demokrati är en process och genom att använda artiklarna i Lomé-konventionen vill vi peka på att förhandlingar kanske , med ett djupt engagemang från de europeiska länderna , kan leda till önskat resultat .
Man skulle också ha kunnat välja att omedelbart avstänga landet från Lomé-biståndet .
Jag tror emellertid att det förfarande som valts ger en del möjligheter på villkor att vi är mycket väl medvetna om vart vi vill komma och att vi även är beredda att ge det här landet effektiv hjälp .
Herr talman , mina kära kolleger !
Den 24 december avbröt en militärstatskupp brutalt demokratin i Elfenbenskusten .
Allt har sagts , nästan allt , om den föregående regimens brister av de talare som har föregått mig .
Anklagelser om korruption har lagts fram .
Det fanns förvisso vissa risker för manipulering av det presidentval som skulle äga rum inom kort .
Jag passar förresten på tillfället att uppmärksamma kammaren på fallet med ett annat land om vilket det inte talas så mycket , Senegal , där ett presidentval kommer att äga rum , som uppvisar samma risker för manipulering som Elfenbenskusten .
Men vi måste vara tydliga .
I Elfenbenskusten liksom på andra ställen kan inte dessa risker vara en ursäkt för det som har hänt där borta .
En statskupp är visserligen inte , och kommer aldrig att vara det , en vinstlott för demokratin .
Mina damer och herrar , parlamentet bör fördöma militärkuppen men det räcker naturligtvis inte .
En övergångsregering har bildats och Europaparlamentet bör göra påtryckningar så att fria och öppna val ordnas redan i juni 2000 , såsom redan begärts av Västafrikas ekonomiska gemenskap , med närvaro av observatörer från världssamfundet och på grundval av trovärdiga vallistor .
Parallellt ber jag att de politiska ledare som arresterades vid statskuppen frisläpps .
Yttrandefrihet och iakttagande av mänskliga rättigheter bör på nytt säkras .
Parlamentet bör under dessa förhållanden nära följa kommissionens åtgärd att begära att samråd inleds om ett eventuellt uppskjutande av samarbetet mellan Europeiska unionen och Elfenbenskusten .
Mina damer och herrar , herr talman , mina kära kolleger , ett återställande av demokrati i Elfenbenskusten bör från och med i dag vara en oförtruten angelägenhet för parlamentet och bortom detta för alla personer som önskar att rätt går före makt .
Herr talman , herr kommissionär !
Demokratin är något mycket skört i Afrika .
Det har ytterligare en gång visat sig i Elfenbenskusten , ett land som ändå var känt som en modell av relativ politisk och ekonomisk stabilitet .
Det är rätt , Bedié-regimen gled snabbt utför mot slutet .
Internationella valutafonden ( IMF ) , Europeiska unionens världsbank , upphävde förra året sitt bistånd till Elfenbenskusten på grund av bristande insyn och öppenhet samt missbruk av statliga medel .
Politiskt gick det också fel .
Presidenten började visa auktoritära och repressiva drag , främst när han likviderade sin viktigaste rival Watara på ett mycket omstritt sätt .
Men är allt det något som berättigar en statskupp ?
Det är nyckelfrågan .
Jag kan inte bli kvitt intrycket att Europeiska unionen intar en mycket mildare hållning gentemot Elfenbenskusten än i andra liknande situationer .
Det är väl ändå svårt att straffa en statskupp i Burundi genom att stödja ett embargo och samtidigt i Elfenbenskusten snabbt övergå till dagordningen .
Genom att inte otvetydigt fördöma denna coup , riskerar man att ge de militära ledarna i Afrika ett alibi för att gripa makten med hjälp av vapen .
Därför måste Europeiska unionen hålla locket på och kräva ett återinförande av rättsstaten och demokratin med hjälp av fria och rättvisa val som conditio sine qua non för varje vidare samarbete med Elfenbenskusten .
Låt oss framför allt inte hantera två olika vikter .
Vad mig anbelangar , herr talman , så finns det inga bra eller dåliga statskupper .
Militära lösningar är definitionsmässigt kortsiktiga lösningar , var i världen de än förekommer . .
( FR ) Herr talman !
Kommissionen , ordförandeskapet och medlemsstaterna har uttryckt sin djupa oro för den upplösning av de offentliga och rättsliga institutionerna som följde på den militära statskuppen .
Europeiska unionen följde redan med särskild uppmärksamhet situationens utveckling i Elfenbenskusten med tanke på arresteringen och fängslandet av oppositionsledarna , den arresteringsorder som utfärdats mot Ouattara , utvecklingen av etniska spänningar samt försämringen av den ekonomiska situationen .
Vårt främsta mål är nu att uppmuntra till ett snabbt återupprättande av rättsstaten och normalt fungerande demokratiska institutioner .
Kommissionen har därför beslutat att inleda det samrådsförfarande som anges i artikel 366b i Lomékonventionen .
Förfarandet är detsamma som det som tillämpades förra året när det gäller Niger och Guinea-Bissau .
Rådet har godkänt förslaget .
Kommissionen och rådet har sänt en inbjudan till Elfenbenskusten .
Elfenbenskustens myndigheter har en frist på fjorton dagar för att besvara inbjudan .
Efteråt bör samrådsförfarandet avslutas inom en månad .
Europaparlamentet kommer att hållas informerat om samrådens förlopp .
Syftena med samråden är följande : att göra en detaljerad utvärdering av situationen i Elfenbenskusten , att betona den vikt som Europeiska unionen fäster vid att de väsentliga delarna av artikel 5 i Lomékonventionen följs , det vill säga respekt för rättsstaten , demokrati och mänskliga rättigheter , att detaljerat känna till Elfenbenskustens avsikter för att säkra respekt för dessa väsentliga faktorer samt nå ett avtal om de åtgärder som kommer att vidtas för att avhjälpa brott mot dessa väsentliga delar .
Kommissionen och rådet arbetar med att förbereda samråden , men jag kan redan säga er att vårt mål är att få ett fast åtagande från Elfenbenskustens myndigheter om återgång till konstitutionell ordning och meddelande om en tidsplan för denna övergång .
Om resultatet av samråden ändå inte är tillfredsställande har Europeiska unionen vid den tidpunkten möjlighet att vidta lämpliga åtgärder , inbegripet ett fullständigt eller partiellt uppskjutande av samarbetet med landet vid behov .
Hittills har inte ett uppskjutande föreslagits eftersom vi vill undvika att bestraffa befolkningarna .
Kort sagt , för närvarande kommer inte något nytt beslut om finansiering att godkännas med undantag av projekt för humanitär hjälp till de minst gynnade befolkningarna .
Avslutningsvis kan jag försäkra er att kommissionen fäster mycket stor vikt vid samråden som kommer att inledas med Elfenbenskusten inom de närmaste dagarna .
Den kommer att uppmärksamt följa situationens utveckling i landet och se till att mänskliga rättigheter respekteras och Europaparlamentet kommer att informeras .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum kl .
17.30 .
 
Mänskliga rättigheter Nästa punkt på dagordningen är gemensam debatt om följande resolutionsförslag : Egypten ( B5-0052 / 2000 ) av Karamanou för PSE-gruppen om det sekteristiska våldet mellan kopter och muslimer i Egypten , ( B5-0056 / 2000 ) av Le Pen m.fl. för TDI-gruppen om massakern på koptiska kristna vid Al-Kochen i Egypten , ( B5-0066 / 2000 ) av Hughes Martin för PPE-DE-gruppen om den senaste tidens religiösa våld i övre Egypten , ( B5-0069 / 2000 ) av Morgantini m.fl. för GUE / NGL-gruppen om den senaste tidens religiösa våld i Egypten , Kina - ( B5-0050 / 2000 ) av Schori och Colom i Naval för PSE-gruppen om Kina , ( B5-0064 / 2000 ) av Haarder m.fl. för ELDR-gruppen om situationen för de mänskliga rättigheterna i Kina , ( B5-0079 / 2000 ) av Gahrton m.fl. för Verts / ALE-gruppen om kränkningar av de mänskliga rättigheterna i Kina , ( B5-0083 / 2000 ) av Van Orden m.fl. för PPE-DE-gruppen om mänskliga rättigheter i Kina , Irak- ( B5-0038 / 2000 ) av Collins för UEN-gruppen om Kuwaitier som hålls fångna i Irak , ( B5-0053 / 2000 ) av Sakellariou för PSE-gruppen om fångar efter kriget i Persiska viken , ( B5-0062 / 2000 ) av Haarder för ELDR-gruppen om fångar i Irak efter krigen i Persiska viken , ( B5-0070 / 2000 ) av Marset Campos m.fl. för GUE / NGL-gruppen om krigsfångar av kuwaitiskt ursprung i Irak , ( B5-0074 / 2000 ) av Boumédiene-Thiery m.fl. för Verts / ALE-gruppen om fångar efter kriget Gulfkriget , ( B5-0084 / 2000 ) av Salafranca Sánchez-Neyra och Grossetête för PPE-DE-gruppen om fångar i Irak efter Gulfkriget , Tchad- ( B5-0078 / 2000 ) av Lannoye m.fl. för Verts / ALE-gruppen om kränkningar av de mänskliga rättigheterna som har samband med oljeutvinnings- och oljeledningsprojektet mellan Tchad och Kamerun , ( B5-0081 / 2000 ) av Howitt och Kinnock för PSE-gruppen om kränkningar av de mänskliga rättigheterna som har samband med olje- och oljeledningsprojektet mellan Tchad och Kamerun , ( B5-0088 / 2000 ) av Novelli för PPE-DE-gruppen om situationen för de mänskliga rättigheterna i Tchad .
Egypten Herr talman !
Med dagens resolution vill jag ge uttryck för den socialistiska gruppens oro för omfattningen av våldet och de blodiga sammanstötningarna mellan anhängare av olika religiösa trossatser .
I Egypten , Indonesien , Nigeria , Libanon , Tjetjenien , Kosovo sätter det religiösa hatet och den religiösa lidelsen själva freden , stabiliteten och utvecklingen på spel .
Millennieskiftet kännetecknades inte bara av fest och firande , utan tyvärr även av blodsoffer - de värsta under senare år - på altaret för det blinda hat som är ett barn av den religiösa fanatismen .
Naturligtvis värdesätter vi den egyptiska regeringens ansträngningar att bemöta extremisterna och hjälpa offren för våldshandlingarna .
Dessa ansträngningar måste emellertid intensifieras , det måste göras en ingående undersökning , de skyldiga måste straffas , och det måste , framför allt , vidtas åtgärder som stärker demokratin , respekten för de mänskliga rättigheterna och toleransen för olika religiösa trossatser .
Ett steg i linje med respekten för de mänskliga rättigheterna skulle naturligtvis vara att avskaffa den medeltida straffmetod som fortfarande tillämpas i Egypten , dödsstraffet .
Vi vet att den egyptiska polisen i början av det nya året med svårighet lyckades få stopp på sammanstötningar i landets södra delar mellan kristna och muslimer , sammanstötningar som kostade 25 människor livet , medan tiotals hus och affärslokaler sattes i brand .
Dessa våldsamheter i Egypten får naturligtvis läggas till tidigare episoder och till fundamentalistiska muslimers blodiga attacker på kristna 1992 och 1997 , som drabbade turismen i Egypten hårt , med negativa följder för landets ekonomiska och sociala utveckling .
Avslutningsvis , med denna resolution skulle jag vilja uppmana rådet och kommissionen att , inom ramen för Meda-programmet , planera för medvetandegörande åtgärder som främjar respekten för de mänskliga rättigheterna och den religiösa toleransen .
Herr talman !
Jag vill först och främst betona att för vår grupp är den brådskande resolutionen framför allt ett starkt påtryckningsmedel för att klara av ett aktuellt problem , där frånvaron av kontroll på politisk nivå kan förstärka en befintlig risk .
I detta fall tror vi dock att den föreslagna texten inte uppfyller kravet på användning av ett brådskande förslag .
Vi förstärks i vår tro genom att vi alla vid granskningen av ärendet såg att rapporterade fakta inte har den politiska omfattning som uttrycks i de första ingresserna i den resolution som man föreslår oss .
Det handlar mer om konflikter av allmän lag i en del av Egypten än om handlingar beroende på religiös antagonism .
Jag måste för övrigt nämna den brist på elegans som det innebär att helt enkelt kopiera ett antal punkter från den skrivelse som hade sänts av talmannen i det egyptiska parlamentet till talmannen i Europaparlamentet .
Att på detta sätt ta över argument som lagts fram av andra för att försvara sig , verkar inte kunna rekommenderas , inte ens intellektuellt .
Eftersom jag dessutom känner till den aggressiva tolkning , som vissa islamistiska miljöer gör av våra initiativ , fruktar vi att i praktiken ge dem ett vapen för att bevisa att Europaparlamentet går för långt i förhållande till en situation som inte berättigar en sådan iver och en sådan politisk beslutsamhet .
Den liberala gruppen kommer därmed inte att rösta för resolutionen .
Vi kommer att lägga ner vår röst samtidigt som vi förbehåller oss rätten att inge ett resolutionsförslag som borde leda till att Europaparlamentet blir litet mindre inskränkt och ser på annat sätt vad som utspelar sig i Egypten och i Nordafrika i sin helhet när det gäller skydd av minoriteters rättigheter och demokratiska rättigheter .
Herr talman , mina kära kolleger !
Ni har framför er ett gemensamt resolutionsförslag rörande de våldsamheter som nyligen försiggått i övre Egypten , i vilka mer än tjugo egyptiska medborgare har dött .
Kära kolleger , ni vet kanske att jag också är föredragande av associeringsavtalet mellan Europeiska unionen och Egypten .
Förhandlingarna om de tekniska ärendena avslutades i juni och vi borde mycket snart få den slutliga texten framlagd .
Avtalet kommer , hoppas jag , att markera tillkomsten av allt närmare förbindelser mellan Egypten , en väsentlig aktör i Mellanöstern och Medelhavsområdet , och unionen .
Den politiska situationen är för närvarande i en gynnsam fas i Mellanöstern och jag ville betona dessa faktorer för att ställa vårt tillvägagångssätt i ett bredare sammanhang .
Med resolutionen vill parlamentet uttrycka sin rörelse inför de händelser som ägt rum men också påminna om att det kommer att vara mycket vaksamt när det gäller mänskliga rättigheter inom ramen för förhandlingarna med våra Medelhavspartner , liksom vi är det med samtliga våra partner .
Vi har placerat skydd av mänskliga rättigheter och demokrati i centrum av vår verksamhet och det är absolut nödvändigt , tror jag , att visa att vi kommer att vara omedgörliga i dessa frågor genom att uppmuntra dem som slår in på den vägen .
Det har inte undgått samtliga kolleger att de egyptiska myndigheterna har reagerat snabbt , som de borde , med att leda en undersökning på platsen och framför allt ordna hjälp till offren för dessa våldsamheter .
President Mubarak ingrep själv mitt uppe i krisen .
Enligt min åsikt är det således tydligt och klart att resolutionen skall ses som ett positivt och uppmuntrande tecken från vår sida , och jag ber samtliga kolleger att godkänna denna text som är resultatet av en kompromiss .
Jag skulle i det avseendet vilja tacka de kolleger som är medundertecknare av förslaget för den goda vilja som de har visat för att komma fram till en gemensam text .
Herr talman , jag skulle vilja avsluta med att säga att texten förvisso har förändrats , och dessutom i förbindelse med de egyptiska myndigheterna , vilket är ett mycket gott tecken .
Herr talman , kära kolleger !
En våg av våldsamheter går fram över Egypten sedan ett tiotal åt tillbaka .
Vi kan dock bara notera den långa tystnaden från såväl världssamfundet som vår europeiska institution .
Egypten spelade visserligen en grundläggande roll i fredsprocessen i Mellanöstern och dess geopolitiska situation gör att ingen egentligen vågar tala om saker som kan framkalla ilska .
Vi kan slutligen bara glädjas åt att en debatt om landet äger rum inom partnerskapet EU-Medelhavsområdet .
Det är däremot beklagligt att det sker av så olyckliga aktuella orsaker .
Vi stöder naturligtvis den egyptiska regeringens ansträngningar i kampen mot den religiösa integrismens uppgång , men denna kamp mot extremism kan inte berättiga ett brott mot det egyptiska folket , i synnerhet av politiska rättigheter .
Den kan inte dölja brotten mot yttrandefrihet och de grundläggande rättigheter som mänskliga rättigheter utgör .
Vi fördömer därför vidmakthållandet av dödsstraff i landet .
Vi ber avslutningsvis rådet att inom ramen för Meda-programmet planera speciella åtgärder för socioekonomisk utveckling , demokratiutveckling och främjande av tolerans mellan samtliga etniska och kulturella minoriteter som utgör det egyptiska samhällets rikedom .
Kina Herr talman !
Det är inte mer än rätt och riktigt att Europaparlamentet för sin oro för situationen för de mänskliga rättigheterna i Kina till protokollet .
Det har varit allt för många fall av religiös intolerans , diskriminering av etniska minoritetsgrupper och fortsatt användning av dödsstraffet för att vi skall kunna ignorera dem .
Vi oroar oss även för de politiska friheterna i Hong Kong och i framtiden i Macao .
Vi gör rätt som sätter press på Kina att förbättra sina meriter .
Det är viktigt att vi i EU fortsätter att göra det .
Jag har dock två kommentarer .
För det första , vi måste akta oss för att i onödan äventyra Kinas anslutning till Världshandelsorganisationen ( WTO ) , eftersom ett WTO-medlemskap på medellång sikt skulle göra mer för att förändra Kinas ekonomi och situationen för de mänskliga rättigheterna i Kina än någonting annat .
Om Kina öppnas upp och integreras i den globala ekonomin , måste det få positiva konsekvenser för de mänskliga rättigheterna .
Många i Kinas ledning känner till och välkomnar detta .
Vi måste vara försiktiga så att vi i våra ansträngningar att nå det bästa inte kastar ut barnet med badvattnet och i slutändan tar ställning för det sämre alternativet .
För det andra , vi måste fortsätta att kritisera Kina .
Jag kommer att fortsätta med det , när så är nödvändigt , men jag hoppas att vi inte kommer att fokusera allt för mycket på Kina , så att vi glömmer bort andra regimer i världen , vars meriter många gånger är lika dåliga , om inte sämre , blir lidande .
Det skulle bara ge Kina en ursäkt att ignorera våra krav .
Herr talman !
Det mest oroande med situationen i Kina är att situationen för de mänskliga rättigheterna i landet , enligt många rapporter , fortsätter att försämras , trots all den dialog som vi har fört med Kina .
Förföljelserna av oliktänkande , arbetsrättsaktivister , religiösa grupper fortsätter , och under de senaste månaderna har vi sett många ledare av Falun Gong-rörelsen interneras utan rättegång .
Det finns ett reellt problem i Kina med tortyr och arbetsläger .
Men , det kanske allvarligaste av allt är att det finns mer än 60 olika brott , av vilka många är icke-våldsbrott , som bestraffas med döden .
Det är de lagliga avrättningarna som är den kanske största anledningen till oro .
1998 registrerade Amnesty International 2 700 dödsdomar och 1 769 bekräftade avrättningar .
Detta är ett mycket allvarligt problem .
Vi måste fortsätta dialogen med Kina ; vi måste anstränga oss för att genom dialog och genom handel öppna upp det kinesiska samhället för västerländska idéer och försöka övertyga dem om det felaktiga i deras metoder .
Herr talman !
Situationen med de mänskliga rättigheterna i Kina har verkligen klart blivit ännu sämre .
Hongkong är ett kapitel för sig som också har ett särskilt " symptomvärde " .
Karmapa Lamas flykt har för sin del kastat ljus över den hårdnande religionsförföljelsen i Kina .
Under dessa förhållanden säger jag ja till Kinas medlemskap i WTO , men hand i hand med detta måste man kräva en ratificering av FN : s konvention om medborgerliga och politiska rättigheter .
Det är viktigt med en retorisk förbindelse till respekten för mänskliga rättigheter , det är det första steget .
Även andra medel måste användas för att EU skall kunna signalera sin oro , och i synnerhet borde man ställa sig bakom den kritiska resolution som Förenta staterna kommer att ta upp vid det kommande mötet med FN : s kommitté för mänskliga rättigheter .
Herr talman !
I och med Martin Lees , den framstående demokratiska ledaren från Hong Kong , närvaro här i Strasbourg och en hög kinesisk WTO-förhandlingsgrupps ankomst till Bryssel på måndag , är frågan om de mänskliga rättigheterna i Kina åter i högsta grad aktuell .
Då vi för fram denna fråga i förgrunden söker vi inte en konfrontation med Kina , ett land som vi hyser stor respekt för och i många avseenden beundrar .
Det är beklagligt att de enorma ekonomiska framsteg som har gjorts i Kina under de senaste tio åren inte har motsvarats av liknande framsteg vad beträffar politisk och religiös frihet samt rättssäkerhet .
Naturligtvis måste det föras en dialog om dessa frågor , men det måste även leda till ett positivt resultat i form av verkliga och väsentliga reformer .
Det är inte godtagbart att säga att västerländska normer inte är tillämpliga i Kina .
De mänskliga rättigheterna är universella , och i detta avseende skiljer sig inte asiatiska värderingar från våra egna värderingar .
I Hong Kong ser vi en urholkning av svårvunna friheter och garantier .
Men kanske är det ingen överraskning att demonstrationer om Tibet är förbjudna där , när de med nöd och näppe är tillåtna i London , om den kinesiske presidenten är på besök .
På det kinesiska fastlandet borde vi gratulera de senaste årens ledarskap till att ha gjort sig av med kommunismen , men i dess plats har vi sett en korrumperad form av kapitalism utan demokrati växa till sig .
Den kinesiska regeringen måste upphöra med att trakassera och fängsla kristna , som Li Dexian i Guandongprovinsen , och att förtrycka buddister i Tibet och på andra platser .
Jag uppmanar de kinesiska myndigheterna att visa kuraget att tillåta demokrater som Martin Lee att resa fritt på det kinesiska fastlandet .
Vi vill se ett Kina som är en fullt integrerad del av det internationella samfundet , med verklig demokrati och rättssäkerhet .
När kommer Kina att upprätta en demokratitidtabell ?
Kommissionär Busquin !
Fastän jag förstår att de mänskliga rättigheterna och handelsförhandlingarna vanligen hanteras var för sig i Europeiska unionen , skulle jag vilja be kommissionen att se till att de kinesiska WTO-förhandlarna i nästa vecka på ett klart och tydligt sätt uppmärksammas på den oro som finns i denna kammare .
Herr talman !
Europeiska unionen är stolt över sitt rykte som försvarare av de mänskliga rättigheterna .
Tyvärr vägrar enskilda medlemsstater att kritisera Kinas brott mot de mänskliga rättigheterna av rädsla för att det skulle skada deras handelsförbindelser .
Detta politiska spel försvagar EU : s moraliska auktoritet att tala om kränkningar av de mänskliga rättigheterna på andra platser i världen .
Jag är föredragande för Hong Kong i detta parlament , och jag är oroad över den mängd incidenter som har inträffat i den delen av världen som , återigen , tyder på kränkningar av de mänskliga rättigheterna .
Avlägsnandet av Cheug Man-Yee som radio- och TV-chef i Hong Kong var ett direkt angrepp på pressfriheten , och beslutet av Hong Kongs SAR-regering att begära en omtolkning av en impopulärt utslag i en högre domstol nyligen träffar rättsstatsprincipen mitt i hjärtat , när högsta domstolens beslut borde ha godtagits .
Behandlingen av Falun Gong-utövare och vägran att tillåta Hong Kongs lagstiftande råd ( LegCo ) att resa till det kinesiska fastlandet är tydliga tecken på de problem som finns kvar i denna delen av världen , och jag kommer att ta upp dessa frågor i mitt betänkande .
Det är mycket viktigt att EU , både som en institution och genom sina medlemsstater , när det är befogat kritiserar Kinas kränkningar av de mänskliga rättigheterna .
Herr talman !
Människorättsläget i Kina har försämrats avsevärt det senaste året .
Tänk bara på det ökande antalet avrättningar , förbudet mot Falun Gong-rörelsen och förtrycket mot Tibet som illustreras av den fjortonåriga tibetanska Karmapa Lamas flykt till Indien helt nyligen .
För den liberala gruppen är måttet nu rågat .
En dialog mellan EU och Kina om de mänskliga rättigheterna är utmärkt , men om resultaten uteblir så måste åtgärder vidtas .
Nu när USA vill stödja FN-resolution om Kina vid det förestående sammanträdet i Genève så uppmanar jag även rådet att göra samma sak och det i enighet .
Historien har nämligen visat hur skadligt det är om vissa medlemsstater låter sina nationella intressen få företräde .
Nederländerna fick uppleva det för tre år sedan då landet i egenskap av ordförandeland för Europeiska unionen gav sitt stöd till en FN-resolution som inte fick ett enhälligt stöd från de övriga medlemsstaterna .
Ekonomiska sanktioner mot Nederländerna blev följden av det .
Den här resolutionen är lackmusprovet för vår herr GUSP , Solana .
På honom vilar den slutgiltiga uppgiften att ena medlemsstaterna om en enda linje den här gången så att rådet går enat i bräschen för universella mänskliga rättigheter .
Herr talman !
Situationen för mänskliga rättigheter i Kina är fortfarande mycket allvarlig .
De mest grundläggande demokratiska och mänskliga rättigheterna respekteras inte .
Försök att formera politisk opposition bekämpas med fängslanden , horribla straff och förvisningar .
Det finns i dag tusentals politiska fångar i landet .
Försök till oberoende , facklig organisering och facklig kamp för arbetandes rättigheter , som inte kontrolleras av kommunistpartiet , tolereras inte .
Det är beklämmande att se hur en stat som säger sig agera i arbetarklassens intresse förtrycker just denna arbetarklass , när den tar till kamp för sina legitima rättigheter .
Dödsstraff utdöms och verkställs i en skrämmande omfattning .
Religionsfriheten respekteras inte .
Förföljelsen av anhängare av Falun Gong-rörelsen är häpnadsväckande och oförsvarlig .
Flera minoritetsfolk , t.ex. tibetanerna , förtrycks och saknar inte bara demokratiska utan också kulturella rättigheter .
Det finns en rad dokumenterade fall av övergrepp och våld från fängelsepersonal och polis .
Det finns därför en mycket god grund för den kritiska resolution som vi skall rösta igenom om en stund .
Jag kommer självklart att rösta för den .
Det innebär inte att jag tycker att alla delar av texten är perfekta .
Jag tycker till exempel att innehållet i punkt 4 delvis skulle ha uttryckts på ett annat sätt .
Jag skulle också gärna haft en skrivning i resolutionen om bristen på fackliga rättigheter i Kina .
Vi ser ju hur den kinesiska regeringen har reagerat mot de strejker och demonstrationer och försök till facklig organisering som vi har sett uppstå den senaste tiden .
Jag skulle också vilja varna för en utveckling som innebär att man tonar ner kritiken mot bristen på mänskliga rättigheter för att uppnå ekonomiska och handelspolitiska fördelar .
Herr talman !
Måndag eftermiddag , när sammanträdet öppnades , bad jag parlamentet och parlamentets talman att sända ett budskap till Texas guvernör för att stoppa en avrättning som skulle äga rum om några dagar .
Mot den bakgrunden är det desto viktigare och skälen desto starkare för att parlamentet i dag skall ägna sig åt situationen i Kina där kränkningen av de mänskliga rättigheterna når sådana enorma proportioner .
Allt detta har redan sagts av mina kolleger och jag kan bara instämma i vad de sagt .
Verkligheten är den att i Kina försämras situationen när det gäller de mänskliga rättigheterna .
Samtidigt som man genomför en besvärlig öppning mot nya ekonomiska system kan vi bevittna en dramatisk försämring när det gäller de mänskliga rättigheterna .
En uppgift från Amnesty International nämner cirka 700 dödsdomar .
En annan siffra från andra källor anger i stället att hela 1 400 dödsdomar verkställdes under förra året .
Oavsett vilken siffra som är den rätta så är det uppenbart att vi står inför något dramatiskt .
Problemet blir då hur man skall kunna hantera detta faktum i unionen och i parlamentet .
Det första vi måste göra , enligt min mening , är att koncentrera oss på nästa session med FN : s kommission för mänskliga rättigheter , den som inleds i Genève den 20 mars med just denna fråga på dagordningen .
Jag frågar mig , och jag frågar denna församling , om man inte kunde begära att unionen , eller till och med parlamentet , fick närvara vid den sessionen .
Men framför allt - och detta har redan sagts - är det inte bara viktigt att unionen gör sin röst hörd utan att den lyckas framföra en gemensam , kraftfull och beslutsam ståndpunkt från de olika medlemsstaterna .
Det är riktigt som redan har sagts : unionens storslagna resolutioner försvagas om de enskilda staterna , av ekonomiska eller kommersiella skäl , handlar tvärtemot .
I det sammanhanget måste vi diskutera en fråga : Kinas ansökan om medlemskap i Världshandelsorganisationen ( WTO ) som , det inser jag , har positiva inslag och som indirekt skulle kunna medföra fördelar , men som också den bör kopplas till en allmän ståndpunkt från FN : s sida och , när det gäller den frågan , en kraftfull uppmaning till Kina att göra framsteg .
I så fall skulle vi kanske kunna gå från uppmaningar , som i och för sig är nödvändiga om än inte tillräckliga , till konkreta handlingar .
Herr talman , herr kommissionär , kära kolleger !
Jag har goda nyheter till er .
Tendensen från de västerländska företagen , således inbegripet de europeiska företagen , att minska investeringarna i Kina betonas och ökar .
Parlamentet är således inte längre ensamt om att opponera sig mot rådet och kommissionen , det råd och den kommission som i åratal har fört en kortsynt politik gentemot Folkrepubliken Kina , en politik grundad liksom i fallet med Sovjetunionen , på samförstånd med en diktaturregim och en kommunistisk regim .
En god nyhet således , vi har allierade : europeiska småföretagare och industrimän .
Vi bör således arbeta för att stärka denna allians och för att äntligen få rådet och kommissionen att inta en sträng och fast ståndpunkt gentemot Folkrepubliken Kina .
Vi måste också ta itu med att skapa ett alternativ eftersom , såsom ni vet , kommunisterna bara förstår maktspråk .
Det är således viktigt att de vet att våra ord kommer att följas av handling och att vår politik kommer att vara trovärdig .
Vi har - och jag tror att vi bör tacka det portugisiska ordförandeskapet - en möjlighet till ett enormt och genomförbart alternativ : Vi kan skapa en strategisk allians med den största och den mest befolkade demokratin i världen Jag talar om Indien och det portugisiska ordförandeskapet , som har tillkännagett att ett första toppmöte EU-Indien skall hållas , ger oss tillfälle att konkret arbeta med att utveckla detta alternativ .
Jag tror att det är det enda initiativ som kan få de kinesiska kommunistiska myndigheterna att förstå att vi inte talar förgäves och att vi allvarligt arbetar för att det kinesiska kommunistväldet äntligen skall störta samman samt att det äntligen skall bli demokrati i Tibet , i Östturkestan , i nedre Mongoliet , som också liksom Tjetjenien är områden som ännu är underkastade en hänsynslös kolonialisering .
Krigsfångar från Gulfkriget i Irak Herr talman !
I dag debatterar vi olika aspekter av den dramatiska frågan om mänskliga rättigheter , och även om vi befinner oss på andra sidan jordklotet så är det nödvändigt att parlamentet låter göra sin röst hörd i ett läge när situationen i Irak fortsätter att vara allvarlig .
Detta land utgör framför allt ett hot för hela regionen och dessutom pågår i Irak en uppenbar kränkning av de mänskliga rättigheterna .
Det är nödvändigt att kräva att de kuwaitiska krigsfångarna släpps fria - enligt de uppgifter som står att få finns det cirka sex hundra krigsfångar som verkar behandlas klart omänskligt - enligt de respektabla röster som hörs i den arabiska världen , som till exempel Arabförbundets generalsekreterare Abdel Meguid , som kräver respekt för mänskliga rättigheter och en förlikning mellan de olika arabstaterna .
Vi får inte glömma att allt detta är följden av den uppenbara kränkning av den nationella suveräniteten som skedde i samband med Iraks aggression mot Kuwait .
I den frågan uppmanar jag Europaparlamentet att göra sin röst hörd och att samtidigt tänka på att det enligt pålitliga källor dessvärre även i Kuwait fortfarande hålls - och det är inte så få - irakiska krigsfångar och att situationen även i det fallet är oroande när det gäller fångarnas mänskliga rättigheter .
Vi måste övertyga Kuwait om att deras krav på att landets rättigheter skall beaktas får mycket större tyngd om landet först uppfyller sina skyldigheter mot humanitetens krav .
Herr talman !
Fallet med de kuwaitiska krigsfångarna är dramatiskt .
De är mer än 600 män och kvinnor som med våld fördes ut ur sitt land av de irakiska styrkorna , när de efter att ha invaderat och ödelagt Kuwait för tio år sedan besegrade lämnade landet .
Det är personer som mycket lätt kan identifieras tack vare en särskild omständighet : Cirka 4 000 fångar fanns instängda i Basra i krigets slutskede .
På en första expedition tog den irakiska militären med sig en del av fångarna , förmodligen till Bagdad .
Just då utbröt det shiitiska upproret i Basra , vilket grymt undertrycktes men som tillät de 3 000 fångar som var kvar att fly och återvända till sitt land .
De som återvände kunde därmed med stor precision fastställa vem som hade varit tillsammans med dem i fångenskap .
Mer än 600 försvunna av en befolkningsmängd på 700 000 är en mycket hög siffra , så pass hög att det har blivit en verklig nationell katastrof .
Trots Röda korsets och Förenta nationernas bemödanden vägrar fortfarande den irakiska regimen att lämna någon som helst information om vad som har hänt dessa människor .
Må vara att de materiella svårigheterna har bemötts av de kuwaitiska myndigheterna , men den mänskliga tragedin är enorm .
Jag har talat med fäder som sett fyra av sina barn försvinna , med kvinnor som såg hur deras män fördes bort och med ungdomar som bara var barn när deras föräldrar anhölls .
Till offrens lidande kan man därför tillägga deras familjers lidande och allvarliga juridiska problem , som till exempel kvinnorna som efter så lång tid inte vet om de är gifta eller änkor .
Min övertygelse är att det internationella samfundet skall kräva ett svar av Irak .
Hur hemskt svaret än är så blir familjernas lidande mindre förskräckligt än den nuvarande ovissheten , outhärdlig för dem och oacceptabel för oss .
Avslutningsvis vill jag insistera på en punkt som tas upp i resolutionsförslaget .
Parlamentet kommer att rekommendera Europeiska unionen och medlemsstaterna att stå fast vid att man innan förbindelserna med Irak normaliseras skall få ett svar av landets regim på frågan om de kuwaitiska krigsfångarna .
För Europeiska socialdemokratiska partiets grupp är detta krav inte mindre viktigt än kravet att Irak skall avväpna sina kärn- , kemiska- och biologiska vapen .
Måtte vår resolution inge hopp för dem som förhoppningsfullt och under förtryck väntar i Kuwait och måtte de som är ansvariga för denna allvarliga situation varnas . )
Herr talman !
I kraft av att kontinuerligt ha motsatt oss alla former av embargon , eftersom det är befolkningen som får lida , men även i kraft av att alltid ha tagit den internationella legaliteten i försvar som en norm för samlevnad och en fredlig lösning av konflikter , kräver vår grupp inte bara att få klarhet i vad som hänt dessa fångar som på ett illegalt sätt tillfångatagits under invasionen av Kuwait , utan också att de förs tillbaka till sitt land - Kuwait - eftersom det är ett sätt att överbrygga övriga problem .
Det är dock inte bara detta det är fråga om - vilket vår kollega Martínez Martínez mycket korrekt beskrev - utan i Irak kränks de mänskliga rättigheterna ideligen , vilket gör det dagliga livet outhärdligt .
Vi menar därför att det passar sig att sätta in den här frågan i ett större sammanhang där Irak måste uppfylla alla villkor som åläggs dem av FN , så att embargot kan hävas och demokratin återinföras .
Herr talman !
Problemet med krigsfångar och försvunna är en del av den katastrofala situationen för de mänskliga och medborgerliga rättigheterna i Irak .
Redan 1992 konstaterade den specielle observatören för FN : s kommitté för mänskliga rättigheter , Max van der Stoel , att Iraks kränkningar av de mänskliga rättigheterna är så allvarliga att de saknar motstycke i världen efter det andra världskriget .
I sin färskaste rapport från förra året tvingas han konstatera att situationen förvärrats ytterligare .
Vi måste ta itu med det här på något sätt .
Krigsfångarna är ett första steg , men förhållandena för allmänheten blir eländigare och vapenkontrollen måste till exempel komma på rätt köl .
Det här fallet med Ekéus , - bråket om det - är ett bra exempel .
Dessa frågor måste man nu ta upp systematiskt .
Herr talman , mina kära kolleger , låt mig sälla mig till de kolleger som redan uttalat sig i debatten för att betona hur outhärdligt problemet är när det gäller familjernas osäkerhet om de sexhundrafem fångarnas och försvunnas öde med hänsyn till mänskliga rättigheter naturligtvis men också individens rätt till värdighet .
Är denna fråga så brännande att det berättigar till en brådskande behandling ?
Ja , enligt min åsikt .
Det är visserligen sant att problemet har funnits där sedan krigsslutet , i mer än nio år , och att de enträgna uppmaningar som vi , parlamentet och Internationella Röda korset har gjort , hittills inte har tillfredsställts .
Jag skulle här vilja godkänna och betona det som vår kollega Martinez just sade .
Vi bör nu ta tillfället i akt för att återuppta förhandlingarna mellan Europeiska unionen och Irak i syfte att eventuellt häva embargot .
Detta tillfälle berättigar i mina ögon att ämnet har förts in för brådskande behandling och det resolutionsförslag som lagts fram för parlamentet för omröstning .
Om vi inte passar på detta tillfälle , tror jag att vi skulle svika vår plikt .
Herr talman !
Den arabiska världen är stadd i rörelse .
Konflikterna i Egypten , vilka vi tidigare har behandlat , har i första hand ingen religiös utan en ekonomisk bakgrund , och den egyptiska staten och de religiösa samfunden anstränger sig ansvarskännande nog för att mildra problemen .
Egypten och Libyen har vad gäller Sudan tagit initiativ för att skapa fred i området , vilket vi bör ge starkt stöd åt .
Trots ett flertal problem , för Syrien en dialog med Israel .
Endast Irak framhärdar i total orörlighet , och jag anser att detta måste få oss att tänka över vår ställning .
Vi måste bedriva en tydlig människorätts- och nedrustningspolitik , självklart just gentemot Saddam Hussein .
Jag vill dock eftertryckligen uttala mitt stöd för vad Morillon sade : vi behöver nu nya förhandlingar .
Vi behöver nya impulser för att faktiskt nå dithän att människorna får hjälp , att framsteg görs , att vi helt konkret knyter möjliga lättnader till helt konkreta framsteg , ända till att nämna namn på förföljda och anhållna personer .
Det måste äntligen tillkomma ett europeiskt initiativ för att sätta fronten i rörelse även här .
Brott mot mänskliga rättigheter i Tchad och Kamerun i samband med de aktuella planerna på en oljeledning Herr talman !
Egentligen är det ett under att den här rörledningen i dag tas upp till diskussion här i parlamentet eftersom det först så mycket lobbyverksamhet för att förhindra det .
Vi är glada att vi kan diskutera den i dag .
Det är i alla fall en början .
Det handlar ju om en omstridd oljeledning mellan Tchad och Kamerun , två länder med mycket dåligt resultat när det gäller mänskliga rättigheter , bekämpandet av fattigdomen , rättssäkerhet .
Vi minns till exempel på nytt Ogoni-området när vi tänker på vilka skadliga följder anläggandet av en oljeledning kan ha om inte de rätta åtgärderna vidtas och de rätta garantierna ges .
Det är till och med så illa att oljeledningen redan nu kastar sin skugga på framtiden , för den i landet som vågar yttra kritik kastas i Tchad helt enkelt i fängelset .
Om det är på det sättet som miljöprotester behandlas i en rättsstat , redan nu , då måste vi undra vad som skulle hända vid värre skador när en korrumperad regim sitter och profiterar på en sådan oljeledning .
Vi vill därför att Europeiska investeringsbanken inte blint följer det som Världsbanken beslutar .
Världsbanken sysslar nämligen med intensiv lobbyverksamhet för att kunna stödja den här oljeledningen och vi vet att de personer , de enda från civil society , som bjöds in att närvara vid ett protestmöte i Amerika , egentligen var lobbyister .
Vi fruktar alltså i högsta grad att de europeiska ledamöterna i Världsbankens styrelse inte kommer att få tid att exakt förbereda sig på en ståndpunkt i den här frågan eftersom det helt enkelt finns så litet objektiv information att tillgå .
Därför ber jag er , herr kommissionär , att se till att Europeiska investeringsbanken inte bidrar till stödet till den här oljeledningen utan att alla sociala och ekologiska försiktighetsåtgärder verkligen vidtagits .
Herr talman !
Vi gör rätt i att behandla oljeledningsprojektet mellan Tchad och Kamerun , som har planerats under flera år , som ett brådskande ärende i dag , både på grund av att det har rapporterats att Världsbanken kan stå i begrepp att fatta sitt beslut och på grund av stor oro över rapporter om trakasserier och hot mot projektets motståndare .
Jag har träffat företrädare för den tchadiska regeringen , som säger , tvärt emot vad de på den andra sidan kammaren hävdar , att de inte har hotat med att dra tillbaka sin inbjudan till parlamentets delegation till Tchad på grund av att vi håller denna debatt .
De hävdar faktiskt att demokratins principer och de mänskliga rättigheterna nu respekteras i samband med detta projekt och att man arbetar i öppenhet .
Men om så är fallet , varför fortsätter vi att få rapporter om överläggningar under vapenhot ?
Varför hotar en tysk icke-statlig organisation på utvecklingsområdet med att dra sig ur på grund av hot och attacker från den tchadiska militärens sida ?
Varför fick en landsflyktig tchadier boende i N ' Djamena den fjärde januari se sitt hem attackeras av tchadiska soldater ?
Om oljeledningsprojektet kännetecknas av öppenhet , varför ifrågasätts dess ändamålsenlighet så fundamentalt i oberoende undersökningar ?
Till exempel , professor Rosenblum på Harvard ifrågasätter effekten på fattigdomen , professor Downing på Arizonas universitet drar slutsatsen att man inte följer Världsbankens riktlinjer för urbefolkningar , och på universitetet i Warwick i mitt eget land anser man att projektet kommer att leda till en potentiell minskning av nationalinkomsten , om hänsyn tas till potentiellt spill och potentiella läckor .
Europaparlamentet gör rätt i att uttrycka sin oro över en världsbank som fortfarande följer de gamla strategierna med privatiseringar , stora infrastrukturprojekt och massexport av jordbruksprodukter som har fått utstå så mycket kritik .
Vad beträffar oljekompanierna själva , varför vill de se miljöskyddskraven lyftas och utvecklingskontrollerna åsidosättas , och till vad behöver de den oinskränkta handlingsrätten i händelse av ett civilt nödläge , som efter vad som påstås kommer att ge dem " en in blanko-fullmakt att agera som en paramilitär styrka " ?
Kan Europeiska investeringsbanken verkligen försvara att man ger 8 miljoner euro direkt till Exxon under dessa omständigheter ?
Vi vill inte ha ett nytt Ogoniland i Afrika .
Herr talman , mina damer och herrar !
För att belysa den debatt som upptar oss skulle jag vilja nämna några siffror för er som talar för sig själva .
När det gäller Tchad först och främst .
Det handlar om den femte fattigaste nationen i världen .
Den förväntade livslängden är under femtio år .
Ett barn av fem dör före fem års ålder , mina damer och herrar .
Årsinkomsten per invånare är 180 dollar .
När det gäller Kamerun är det knappast bättre med en inkomst per invånare på omkring 650 dollar .
Varför nämner jag dessa siffror ?
Helt enkelt för att de uttrycker och visar på den absoluta nödvändigheten att ge dessa länder , i synnerhet Tchad , de utvecklingsmöjligheter som de har rätt till .
Jag tror att det är i detta sammanhang som vi noggrant bör granska det stora projektet för exploatering av oljefälten i södra Tchad samt byggandet av en oljeledning mellan Tchad och Kameruns kuster .
Projektet anses för närvarande väsentligt för dessa båda länders utveckling .
Vi kan bara ett ögonblick tänka oss att med det resultat man väntar sig av exploateringen av oljefälten skulle Tchads bruttonationalprodukt kunna öka med nära tio procent och ge vinster åt landet på mellan fem och tio miljarder dollar .
Världsbanken , som ännu inte har avgett sin slutliga åsikt , följer mycket nära projektet och hjälper Tchad med genomförandet .
De tre främsta frågorna , det vill säga miljö , sociala problem och förvaltning av inkomsterna från projektet , är sedan nära fyra år föremål för mycket djupa undersökningar .
Det kan bedömas av följande : 900 sammanträden har hållits om oljeledningens sträckning , 40 000 personer har gett sin åsikt och 250 icke-statliga organisationer har tillfrågats .
Direktören för en av dem , World Wide Fund for Nature ( Världsnaturfonden ) , anger till och med att när det gäller miljö är anläggningsprojektet för oljeledningen ett av de bästa i världen .
Vi måste ändå naturligtvis fortsätta att nära följa projektets konsekvenser och se till att det blir minsta möjliga skador i fråga om miljö och på det mänskliga planet .
Det är skälet för debatten i dag .
Om Världsbanken , vars kritik jag har svårt att förstå , händelsevis efter de kompletterande undersökningarna skulle ge ett avslag , kan det inte bli fråga om att fortsätta .
Om institutionen däremot slutligen stöder programmet kommer det att betyda att våra legitima farhågor kan lätta och det betyder också att utvecklingen av de fattiga länderna , som är föremål för många tal här , för en gångs skull konkret kommer att bli föremål för vår uppmärksamhet .
Mina damer och herrar , mänskliga rättigheter är också rättigheter till utveckling .
Vi har dåliga erfarenheter av oljeprojekt i Afrika .
Därför bör vi mycket kritiskt bedöma den här frågan på grundval av relevans för utvecklingen och miljövillkor .
Den planerade oljeledningen genom Tchad och Kamerun kan skapa viktiga inkomster för de här länderna som inte kan skapas på något annat sätt .
Min grupp konstaterar att det fanns viktiga invändningar mot de ursprungliga planerna .
Planerna har nu anpassats på alla dessa punkter och den stora frågan är om det nu är tillräckligt .
Vi anser att det här projektet på kort sikt kan gå igenom först när det står obestridligt fast att de strängaste kriterier uppfylls och även Världsbanken uttryckligen och otvetydigt har givit sitt godkännande .
Samtidigt måste det stå helt klart att inga mänskliga rättigheter kränks .
Bara om det är fallet får Europeiska investeringsbanken ge sina lån .
För vår grupp är det här ett test case om det också går att få goda erfarenheter av oljeprojekt i Afrika . .
( FR ) Herr talman , kommissionen är orolig för de våldsutbrott , som de kristna befolkningarna i området Al Kocheh i övre Egypten blivit offer för , och beklagar förlusten av ett stort antal människors liv .
Den konstaterar att den egyptiska regeringen redan har vidtagit åtgärder för att återställa lugnet i området och gläder sig åt dess åtagande att ställa de ansvariga inför rätta .
Kommissionen väntar med intresse på den egyptiska åklagarens preliminära rapport som är planerad till nästa vecka .
Enligt de första meddelandena är de senaste händelserna helt olika händelserna från augusti 1998 , som huvudsakligen utlöstes av ordningsstyrkornas våldsamma och inkompetenta reaktion och inte av ett sekteristiskt uppförande från deras sida .
De senaste händelserna verkar däremot ha en religiös prägel , även om de utlöstes av en enkel handelstvist .
I övre Egypten liksom på andra håll kan den kroniska underutvecklingen på ett farligt sätt intensifiera religiösa spänningar och det är därför som de åtgärder som syftar till att återställa lugnet mellan de olika samfunden bör gå hand i hand med den socioekonomiska utvecklingen .
Kommissionen anstränger sig framför allt i sitt samarbete med Egypten att finna en balans mellan åtgärder för ekonomisk modernisering och sociala åtgärder , inbegripet åtgärder för kamp mot fattigdom samt främjande av det civila samhället och mänskliga rättigheter .
Övre Egypten är ett av de områden till vilka de sociala åtgärderna och åtgärderna för kampen mot fattigdomen riktas .
När det gäller Kina delar kommissionen parlamentsledamöternas oro i fråga om situationen för mänskliga rättigheter i Kina och i synnerhet i Tibet .
Dessa frågor togs upp på högsta nivå vid det andra toppmötet EU-Kina den 21 december 1999 i Peking .
Unionen gjorde också den 14 januari en formell uppvaktning av det kinesiska utrikesministeriet och uttryckte sin djupa oro för de politiska dissidenternas öde , religionsfrihet för medlemmar av de kristna kyrkorna och den behandling som ges åt vissa troende från rörelsen Falun Gong .
Dessa frågor liksom fängelsevillkor , arbetsläger , yttrandefrihet , föreningsrätt samt kvinnors och etniska minoriteters rättigheter kommer också att stå på föredragningslistan vid nästa dialogsammanträde EU-Kina om mänskliga rättigheter som kommer att hållas den 25 februari i Lissabon .
Mot bakgrund av resultatet av sammanträdena och dialogen kommer unionen efteråt att ta ståndpunkt inför nästa sammanträde av Förenta nationernas kommission för mänskliga rättigheter .
Unionen anser att en förbättring av situationen för mänskliga rättigheter i Kina samt förhandlingarna om landets anslutning till WTO utgör två stora utmaningar som det är nödvändigt att behandla åtskilt med hjälp av speciella instrument och inom ramen för specifika organisationer .
I allmänhet kan sägas att kommissionen är av den åsikten att en ekonomisk öppning och en liberalisering av handelsutbytet , som skall påskynda Kinas anslutning till WTO , i längden utgör ett positivt underlag för en gynnsam utveckling av mänskliga rättigheter , ett stärkande av det civila samhället och uppbyggnaden av en rättsstat i Kina och den kommer att vara särskilt uppmärksam på de senare aspekterna inom ramen för dialogen med WTO .
Frågan om Tibet har redan i stort tagits upp med de kinesiska myndigheterna via de nu befintliga kommunikationskanalerna .
Trojkans ambassadörer gjorde för övrigt en observationsresa till Tibet 1998 och kommissionen åtar sig att fortsätta på den vägen .
När det gäller problemet med krigsfångarna från Gulfkriget i Irak oroar sig kommissionen på samma sätt som parlamentet för bristen på samarbete från Iraks sida i ärendet om de försvunna från Kuwait och bedömer de outhärdliga effekterna av situationen för familjerna .
Kommissionen anmodar Irak att respektera resolutionerna av FN : s säkerhetsråd i frågan och , såsom ni betonade , har Internationella Rödakorskommittén fått ansvaret för ärendet om de försvunna från Kuweit , i enlighet , med FN : s resolutioner .
Men Irak vägrar tyvärr att samarbeta , till och med genom denna internationella organisation .
Kommissionen stöder Internationella Rödakorskommitténs ansträngningar och eftersom kommissionen inte har avtalsenliga förbindelser med Irak , finns det således inte någon officiell dialog med den irakiska regeringen .
Dessutom skulle jag vilja försäkra er om att kommissionen helt och fullt instämmer med de sanktioner som införts av Förenta nationerna och som utgör ett svar på den dramatiska situationen för mänskliga rättigheter i landet .
Men såsom vissa av er har betonat , och där tror jag också att vi har en viktig punkt , trots Iraks överträdelser av FN : s säkerhetsråds resolutioner kommer kommissionen att fortsätta att genom ECHO ge humanitär hjälp till irakierna för att lätta deras lidanden .
Kommissionen är den främsta givaren av humanitär hjälp till Irak med ett belopp på 240 miljoner euro sedan 1991 och inom ramen för programmet för år 2000 har ECHO avsatt tio miljoner euro för humanitär hjälp till Irak .
Vi gör således en åtskillnad mellan befolkningarna och överträdelserna av mänskliga rättigheter som är Iraks sätt att handla .
Kommissionen kommer att stödja samtliga åtgärder i frågan .
När det slutligen gäller överträdelserna av mänskliga rättigheter i Tchad och Kamerun i samband med de aktuella planerna på en oljeledning , följer Europeiska kommissionen uppmärksamt situationen beträffande fördjupandet av den demokratiska processen , skydd av mänskliga rättigheter samt stärkandet av rättsstaten .
Kommissionen har också uppmärksamheten på det planerade projektet för oljeexploatering i södra delen av landet , som kommer att gå igenom Kamerun .
Kommissionen är inte direkt berörd av projektfinansieringen .
Men vid flera tillfällen har den visat sin förståelse för Tchads rätt att exploatera sin enda resurs , förutsatt att nödvändiga försiktighetsåtgärder vidtas i fråga om miljöskydd och skydd av de lokala befolkningarnas rättigheter , å ena sidan , och den verkliga användningen av landets framtida oljeinkomster , å andra sidan .
Vi kommer att se till att dessa betänkligheter vidarebefordras till Europeiska investeringsbanken .
I Tchad kommer oljeexploateringen att kunna bli en viktig faktor för utveckling och stärkande av rättsstaten om dessa inkomster används förnuftigt .
Europeiska kommissionen kommer därför att anstränga sig att uppmuntra regeringen att fortsätta dialogen om de frågor som uppstår i samband med oljeprojektet med de främsta partnerna i landet , inbegripet kommissionen själv , och att nära knyta de lokala myndigheterna och icke-statliga organisationer till de förberedande åtgärderna .
Det bör göras så att de framsteg som redan genomförts i fråga om de mest kritiska punkterna i oljeprojektet i förekommande fall kan stärkas .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum om en stund kl.17.30.
 
Situationen på Moluckerna ( Indonesien ) Nästa punkt på föredragningslistan är debatten om sex resolutionsförslag rörande situationen på Moluckerna .
B5-0034 / 00 av Maij-Weggen för PPE-DE-gruppen om Moluckerna och Indonesien , B5-0054 / 00 av Schori och Wiersma för PSE-gruppen om Moluckerna , B5-0059 / 00 av Maaten för ELDR-gruppen om Moluckerna , B5-0071 / 00 av Vinci och Brie för GUE / NGL-gruppen om situationen på Moluckerna i Indonesien , B5-0073 / 00 av Lagendijk för Verts / ALE-gruppen om Moluckerna , B5-0085 / 00 av Maij-Weggen m.fl. för PPE-DE-gruppen om Moluckerna och Indonesien .
Herr talman !
Det här är faktiskt tredje gången på ett halvår som vi måste fästa komissionens uppmärksamhet på Moluckerna .
Vi är missnöjda med komissionens hittills mycket begränsade reaktioner .
Våldsamheterna på Moluckerna började redan förra året .
Inledningsvis stod de i skuggan av det som hände i Östtimor men det gör inte situationen på Moluckerna mindre allvarlig .
I oktober talade vi om hundratals döda .
Nu , tre månader senare , är det tal om tusentals döda och ännu fler skadade och flyktingar .
Naturligtvis är orsakerna av olika art .
Området har blivit ekonomiskt försummat under Suhartus regim och den regimen har också bidragit till att en betänklig migrationspolitik förs .
Det som emellertid är allvarligare är att det nu finns provokatörer , precis som i Östtimor , som uppviglar befolkningen mot varandra och att militären , tyvärr , spelar en betänklig roll .
Det senare bekräftades också i går i en intervju med president Wahid på den nederländska televisionen , där han sade att även militären uppvisar ett beteende som är klandervärt .
I vår resolution riktas kritiken med eftertryck inte på den nya regeringen i Indonesien .
Den gör ärligen sitt bästa för att återupprätta demokratin och göra något åt kränkningarna av de mänskliga rättigheterna .
Det onda i Indonesien verkar mer ligga hos aggressiva muslimorganisationer och provokatörer från militären .
Vad kan Europeiska unionen göra ?
Till att börja med skulle den kunna framföra en varning , såsom även Holbrooke har gjort , om att en statskupp av militären i Indonesien inte kommer att tolereras .
För det andra skulle en oberoende undersökningskommission kunna tillsättas och skickas till Indonesien , helst med ett mandat från FN , för att utreda vad som har hänt under de senaste månaderna .
Samtidigt skulle en förlikningskommitté kunna skickas till området för att försona muslimer och kristna med varandra .
President Wahid har redan bett om det och även nämnt ett namn .
Det skulle vara bra om Europeiska unionen stödde ett sådant initiativ .
Det behövs naturligtvis mycket mer hjälp än den som nu ges .
Avslutningsvis skulle jag vilja peka på att vapenembargot måste förlängas .
Det finns det all anledning till så länge militärens roll är så tvivelaktig .
Jag vill påpeka att striderna och våldet på Moluckerna redan har hållit på alldeles för länge .
I Nederländerna finns en stor gemenskap med rötter i Moluckerna .
Det är en europeisk gemenskap och av det skälet kan Europeiska unionen inte blunda för problemen på Moluckerna .
Vi uppmanar rådet och kommissionen att visa mycket mer handlingskraft än de visat hittills .
Herr talman !
Jag talar för min kollega Wiersma .
Herr talman !
Ministerrådets beslut att upphäva vapenembargot mot Indonesien är kortsiktigt och förhastat .
Indonesien har nu tagit sina första steg på väg mot ett demokratiskt samhälle .
Men såsom den amerikanske FN-ambassadören Holbrooke återigen underströk den här veckan med sin varning till den indonesiska militären så är övergången till ett fullvärdigt demokratiskt statsskick ännu inte ett avgjort lopp .
Den roll som den indonesiska militären spelat under oroligheterna i Östtimor har ännu inte klarats ut .
Spänningen ökar i Indonesien .
Jakarta har ingen kontroll över situationen på Moluckerna .
Det klargjorde min kollega Maat alldeles nyss .
Stora grupper medborgare känner sig inte längre trygga .
Med ett för tidigt upphävande av vapenembargot mot Indonesien riskerar Europa att bli medskyldigt till en upptrappning av våldet .
Därför anser vi att rådet bör ompröva sitt beslut .
Vi uppmanar nu verkligen medlemsstaterna att , i väntan på ett nytt beslut , inte återuppta vapenleveranserna .
Vi ber kommissionen och rådet att vidta fyra åtgärder .
För det första bör Europeiska unionen skicka en delegation till Jakarta för att tillsammans med Wahids regering diskutera en utväg ur den här krisen .
För det andra bör EU träffa överenskommelser med den indonesiska regeringen om att tillåta oberoende observatörer på Moluckerna .
För det tredje bör det ges mer humanitär hjälp till alla delar av befolkningen .
Slutligen bör det via FN och de icke-statliga organisationerna skickas mer hjälp till flyktingar och hemlösa .
Får jag avslutningsvis även tala om hur besvikna vi , den nederländska socialdemokratiska delegationen , är över vår utrikesminister som inte vet hur han skall hålla sig i den här debatten .
Först var han för ett vapenembargo men efter ett besök i Jakarta så tog han tillbaka det .
Europeiska unionen måste handla nu innan det blir för sent .
Jag uppmanar särskilt det portugisiska ordförandeskapet i Europeiska unionen att ta initiativet .
Herr talman !
Jag blev mycket arg när jag i måndags hörde att ministerrådet inte kommer att förlänga vapenembargot .
Jag har förstått att Frankrike , Italien , Spanien och Belgien ville att det skulle hävas , och Storbritannien undvek , som vanligt , att ta ställning .
Så mycket var den etiska utrikespolitiken värd .
Men jag uppmanar EU : s ministerråd att tänka om .
Under tiden bör ingen medlemsstat återuppta vapenhandeln .
Det ger fel signal vid fel tidpunkt .
Till och med den indonesiska kabinettministern har sagt att det var fel beslut .
Demokratin är ömtålig .
Hotet om en armékupp finns där , våldet på Moluckerna förvärras , och vi hör nu från Lombok att tolv kyrkor har bränts ned och att 5 000 människor har flytt , och återigen finns det rapporter om att armén har varit inblandad .
Jag vädjar till ministerrådet att återställa vapenembargot för att främja stabiliteten i Indonesien .
Herr talman !
Den nuvarande enhetsstaten Indonesien är en produkt av 350 års nederländsk kolonialmakt .
Den till kristendomen omvända befolkningen på Moluckerna rekryterades till den kolonialarmé som skulle hålla de andra befolkningsgrupperna under nederländsk makt .
För femtio år sedan flyttade en stor del av Sydmoluckernas befolkning till Nederländerna och sedan dess har en stor utvandring skett från det tätbefolkade Java till de övriga öarna .
Det gör att de av Moluckernas befolkning som stannade kvar har blivit en minoritet i sitt eget område .
Den indonesiska militären genomförde år 1965 en statskupp som troligen kostade en miljon människor livet .
Inte heller efter valet 1999 lyder militären under någon demokratisk auktoritet .
Den agerar som anstiftare av motsättningar mellan befolkningsgrupper .
I måndags bad jag rådet behålla vapenembargot mot Indonesien .
Det gör det möjligt för nederländska och franska företag att inte göra sig skyldiga till kontraktsbrott när de inte verkställer tidigare beställningar av militär utrustning .
Europa bör inte förvåna sig över att det utbryter fler inbördeskrig i Indonesien om vi vägrar inse att militären har intresse av att det utkämpas etniska och religiösa konflikter som har sitt ursprung i den koloniala historien .
Herr talman !
Sista gången som vi i den här salen talade om Moluckerna så sade jag att vi just då talade om Moluckerna , men att jag var rädd att vi inom kort skulle behöva diskutera andra delar av Indonesien .
Det var , för tydlighetens skull , inget förnekande av just den diskussionen och de specifika problemen på Moluckerna utan en analys av problemet i Indonesien som sträcker sig mycket längre än endast Moluckerna och som är mycket strukturellt och djupgående .
Tyvärr måste jag säga att jag fick rätt .
I de senaste rapporterna talas det om att avskyvärda scener nu även utspelar sig på Lombok , scener som påminner om Moluckerna och andra platser i Indonesien där strider blossat upp och där nästa oroskälla skall visa sig , till exempel på Sulawesi .
Allt det här är konsekvenser , bland annat av orkestrerade hatkampanjer , bland annat till och med av ordföranden i den lagstiftande församlingen .
Däremot är president Wahids reaktion hoppingivande .
Jag tror också att Europaparlamentet bör stödja honom i kampen mot intolerans och för en återhållsam liberal form av islam men även främst i hans kamp mot stora delar av armén som inte gör tillräckligt mot orosstiftare och som , ännu värre , vägrar ta sitt ansvar , till exempel för sin egen roll i Östtimor .
Vad jag emellertid inte kan inse är att president Wahid bör få stöd genom att man återupptar vapenleveranserna .
EU har diverse möjligheter att påverka processen i Indonesien .
Mina kolleger har redan tagit upp det : observatörer , humanitärt bistånd .
Till det hör dock också , och det är främst en uppmaning till medlemsstaterna , ett vapenembargo .
Det som behövs i Indonesien är att militärens roll tvingas tillbaka .
Den skall inte förstärkas genom leverans av ännu mer vapen .
Herr talman , herr kommissionär , ärade ledamöter !
Jag noterar att Europeiska rådet , när det beslutar att avskaffa vapenembargot mot Indonesien , intar motsatt ståndpunkt mot vad parlamentet mycket enhälligt rekommenderade förra månaden .
Skälen som ledde fram till embargot har inte förändrats , sedan parlamentets ståndpunkt , vi har situationen på Moluckerna , vilket uttrycks bra i den gemensamma resolutionstexten som vi diskuterar .
Som jag för en månad sedan hävdade är den nuvarande indonesiska regeringen , som utsetts i fria val och riktar in sig på de demokratiska värdena , bland vilka jag vill betona respekten för de mänskliga rättigheterna , förtjänt av uppskattning och solidaritet från det internationella samfundet .
Situationen på Moluckerna , som inte är ett isolerat fall i Indonesien och en följd av den migrationspolitik som Suharto bedrev , till vilken de indonesiska väpnade styrkornas nuvarande agerande kan räknas , ett agerande som är en upprepning av det som skedde i Östtimor under den värsta perioden , som om ingenting hade hänt i landet , motiverar en försiktighet och vissa kriterier för hur vi skall uttrycka solidariteten .
Jag stöder alltså det nödvändiga förstärkta internationella samarbetet genom framför allt humanitär hjälp och utvecklingsbidrag till Indonesien , vilket är ett sätt att visa vår positiva värdering av den nuvarande regeringens demokratiska karaktär vilket kan bidra till att öka dess förmåga att hävda sig .
Jag avvisar vapenförsäljning som går till de väpnade styrkorna som ännu inte har förstått sin status i en rättsstat , vilken placerar dem under regeringens överhöghet .
Med tanke på omständigheterna är den säkra signal vi kan ge att bibehålla vapenembargot mot Indonesien .
Det skulle vara katastrofalt om militären återtog makten i Indonesien .
Därför måste Europa stödja president Wahid i hans försök att återskapa freden på Moluckerna .
Hittills har Europeiska unionen kommit till korta i det avseendet .
Vi måste ge mer humanitärt bistånd och hjälpa indoneserna att få muslimer och kristna att sitta ner vid förhandlingsbordet .
En europeisk delegation , till exempel under ledning av Nederländernas före detta premiärminister Lubbers , skulle kunna förrätta ett bra jobb .
ELDR-gruppen beklagar att vapenembargot inte förlängs .
Det är fortfarande fråga om en spänningshärd och om kränkande av de mänskliga rättigheterna .
Rådet ( allmänna frågor ) håller sig alltså inte till de egna europeiska kriterierna för ett vapenembargo .
Europeiska unionens beslut spelar militären i händerna och det ju just det som inte får hända .
Herr talman , herr kommissionär , kära kolleger !
Efter Egypten , Turkiet och Mellanöstern i allmänhet sprider sig nu påtryckningarna , övergreppen och morden på kristna till Asien .
Det är dags att vi med kraft uttrycker vår revolt inför dessa upprörande händelser .
Religionsbudskapet i Bibeln är ändå tydligt , enkelt och positivt .
Det går inte att föreställa sig att det skall snedvridas för att berättiga till sådana fasor .
Islamismen har genom en lång och regelbunden påtryckning redan tvingat de flesta kristna i Orienten till exil .
Vad gör vi konkret för att stödja dem ?
En mängd sammanslutningar i Frankrike och Europa försöker komma dem till hjälp , så att exil inte är den enda lösningen som återstår för dem .
Jag hyllar dem varmt här i dag .
Vilken utarmning och vilken förlust för dessa länder .
De kristna som finns i dessa länder sedan långt före islams utbredning är också deras kulturella rötter .
På Moluckerna är situationen förvisso annorlunda eftersom den indonesiska regeringen utan framgång försöker kontrollera situationen , oförmögen som den uppenbarligen är att kontrollera sina egna väpnade styrkor , och därför är det absolut nödvändigt att inte ta bort vapenembargot .
Man kan frukta att de kristna än en gång kommer att tjäna som syndabock där till priset av sitt liv för kriser som övergår deras förstånd .
Den indonesiska statens kris har djupa ekonomiska , sociala , politiska och religiösa rötter .
Kära kolleger , därmed uttrycker vår grupp med full kraft sin fasa inför allt som försiggår på Moluckerna , liksom den gjorde inför det som hände i Östtimor , och sin djupa oro för det öde som väntar de kristna i Mellanöstern och nu i Asien .
Herr talman !
President Wahid förnekar fortfarande att konflikten på Moluckerna har utmynnat i en kris .
Det religiösa våldet där beror enligt honom på en våldsbenägen minoritet , de så kallade " dark forces " , som ständigt blåser nytt liv i konflikten .
Nya bilder och underrättelser ger annars en annan bild .
Anstiftande av bränder i kyrkor och moskéer i stor skala och upprepade uppmaningar till ett heligt krig , jihad , anger hur allvarligt läget är .
Att våldsamheterna utbrett sig till Lombok och Sulawesi är också mycket oroväckande .
De inbördes blodigheterna på Moluckerna har redan hållit på i ett år nu .
Det är naturligtvis frestande att söka efter de direkt skyldiga till en sådan konflikt .
Den indonesiska pressen håller också på för fullt med det .
Det kan dock ifrågasättas om det verkligen bidrar till en lösning av konflikterna .
Just nu verkar det till och med som om media bara ytterligare uppmuntrar våldet .
Underrättelserna är inte sällan anledning till nya attacker .
Förutom pressen så spelar även militären en tvivelaktig roll .
Både muslimer och kristna kommer med beskyllningar mot militären .
Wahid försöker väl få kontrollen över armén men det har han ännu inte lyckats med helt .
Därför verkar det inte så klokt att nu upphäva vapenembargot mot Indonesien .
I den gemensamma resolutionen uppmanas rådet , kommissionen och parlamentet att via delegationer bidra till en lösning på konflikterna i Indonesien .
Vi kan naturligtvis inte kliva in där och föreskriva ett antal lösningar .
I det indonesiska samhället måste etniska och religiösa minoriteter och alla andra samhällsaktörer ta tag i uppbyggandet av ett civilt samhälle .
Humanitärt bistånd måste erbjudas så snabbt som möjligt . .
( FR ) Herr talman , kommissionen delar den åsikt som uttryckts av parlamentet i resolutionsförslaget .
Både vad som gäller den indonesiska regeringens fasta åtaganden att främja demokrati och respekt för mänskliga rättigheter och nödvändigheten att stödja den indonesiska regeringen i dess ansträngningar att begränsa våldet och återupprätta mänskliga rättigheter i provinsen Moluckerna .
Beträffande den fredliga dialogen såsom instrument för att återställa freden mellan de muslimska och de kristna samfunden är kommissionen övertygad om att den aktuella situationen - som är så oroande - kräver en insats av världssamfundet .
Det är i detta syfte vi måste stödja den indonesiska regeringen och undvika alla typer av straffreaktioner .
Ordförandeskapets senaste förklaring från den 17 januari återspeglar i hög grad denna attityd och på kommissionär Pattens vägnar kan jag försäkra er att kommissionen instämmer med de tankar som uttrycks i förklaringen .
Rådet ( allmänna frågor ) som är planerat till måndagen den 24 januari kommer emellertid att vara rätt tillfälle för att granska parlamentets begäran .
Det kommande besöket av den indonesiska presidenten i Bryssel , liksom i andra europeiska huvudstäder , kommer dessutom att ge tillfälle att försäkra honom och hans regering om vår vilja att sätta in alla nödvändiga ansträngningar för att problemet skall lösas på fredlig väg .
När det gäller humanitär hjälp är ECHO och kommissionen fullt ut beredda på att stärka den .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum kl .
17.30 .
 
Venezuela Nästa punkt på föredragningslistan är debatten om följande sex resolutionsförslag : B5-0047 / 00 av ledamöterna Muscardini och Ribeiro e Castro för UEN-gruppen om Venezuela .
B5-0055 / 00 av Medina Ortega för PSE-gruppen om de katastrofala översvämningarna i Venezuela .
B5-0060 / 00 av ledamöterna Sánchez García och Di Pietro för ELDR-gruppen om de katastrofala översvämningarna i Venezuela .
B5-0072 / 00 av ledamöterna Wurtz med flera för GUE / NGL-gruppen om översvämningarna i Venezuela .
B5-0076 / 00 av Knörr Borràs och Lipietz för Verts / ALE-gruppen om de katastrofala översvämningarna i Venezuela .
B5-0086 / 00 av Marques och Salafranca Sánchez-Neyra för PPE-gruppen om katastrofen i Venezuela .
Herr talman !
Den som följer den brådskande debatten här i parlamentet tycker nog att det ser ut som om Europas historia återupprepas .
Med andra ord fick vi under den föregående debatten höra mycket nederländska och nu fruktar jag att kommissionären kommer att få höra mycket spanska eftersom vi talar om Venezuela .
Det som händer är att Europas historia upprepar sig .
Det vill säga , de européer som åkte ut och ockuperade världen påverkas nu på ett eller annat sätt av det som händer där ute .
När vi talar , även om det i första hand för kommissionären kan verka som en enda lång klagovisa , så talar vi som företrädare för våra väljare .
I mitt land , och i den region jag kommer från - Kanarieöarna - så känns katastrofen i Venezuela som om den inträffat i vårt eget område .
Jag beklagar att Busquin , en storslagen kommissionär och politiker som väl känner till problemen , inte är den kommissionär som ansvarar för ärendet i fråga .
Han hade förmodligen redan hunnit skrivit ned svaret och det jag kommer att säga skulle inte influera honom , det är jag säker på .
Jag hoppas dock att han åtminstone läser igenom förslaget till resolution och tittar på några av de frågor som oroar oss .
Katastrofen i Venezuela är inte en vanlig katastrof .
Vi talar här om 50 000 försvunna - i stort sett 50 000 döda - , ett lands undergång - Vargas land - där Maiquetía flygplats och La Guaira hamn ligger , Venezuelas port eller hall .
Landet måste återuppbyggas och på ett sätt som gör att en katastrof aldrig mer kan inträffa .
Katastrofen inträffade nämligen inte på grund av myndigheters försumlighet .
Den orsakades av en bergstopps ras - bergstoppen i Avila nationalpark - något som måste uppmärksammas vid återuppbyggnaden .
Jag hoppas att kommissionen beaktar parlamentets synpunkter och att man kan beakta möjligheten av att sammankalla en " givarkonferens " , eller något liknande , tillsammans med andra organisationer och länder så att vi kan bistå den venezuelanska regeringen i återuppbyggnaden av en mycket viktig del av landet . )
Herr talman , herr kommissionär , ärade kollegor !
Vi som kommer från Kanarieöarna , en ultraperifer region i Europeiska unionen , berörs väldigt mycket av allt som händer i Venezuela .
I mitten av förra århundradet tvingades nämligen tusentals kanariebor att emigrera dit , så många så att vi faktiskt betraktar Venezuela som vår åttonde ö .
Vi berörs väldigt mycket av den katastrof som inträffade i Vargas och Mirandas land i mitten av december förra året .
En katastrof som förorsakades av störtregn , laviner och översvämningar vid den venezolanska kusten , vid foten av Avila , en nationalpark där jag själv haft glädjen att arbeta .
De mänskliga förlusterna var höga , liksom skadorna , de materiella förlusterna uppgick till tusentals miljoner euro .
Med exemplarisk solidaritet reagerade vi alla inför katastrofens magnitud , från Europa och Amerika skickades humanitärt och ekonomiskt bistånd .
Med andra ord kom den internationella reaktionen snabbt på alla nivåer , inklusive från Europeiska kommissionen , några medlemsstater och några spanska provinser som står särskilt nära Venezuela .
När nu väl inledningsfasen är över , och trots andra naturincidenter de senaste dagarna , är det mer än någonsin nödvändigt att rehabilitera och återuppbygga bostäder , utrustning och berörd infrastruktur - förutom de hydrologiska korrigeringarna - samt att moraliskt och ekonomiskt ge naturkatastrofens offer vårt stöd , det är nämligen en av de största tragedier som inträffat i Latinamerikas historia , särskilt när det gäller Venezuela .
Vi har därför alla lagt fram ett förslag till resolution där vi först och främst från Europeiska unionens sida i samarbete med medlemsstaterna och andra institutioner försöker uppnå en teknisk och finansiell plan , bland annat , för att mildra och kompensera naturkatastrofens effekter .
Jag kan garantera att katastrofen i Venezuela den här gången har blivit en " aktuell , brådskande och synnerligen viktig " fråga . )
Herr talman !
Det tråkiga är att vi de korta stunder vi ses tvingas tala om olika katastrofer som ödelägger vissa delar av världen , en del mer än andra , och kanske också om att länder med stor fattigdom och svag infrastruktur får betala ett högre pris än om de vore starkare .
Detsamma kan sägas om invånarna , i fallet med Venezuela måste man , som i fallet Mitch , tala om de många dödsoffren .
Givetvis uppmanar vi de europeiska institutionerna att bistå ekonomiskt - och de har redan bistått , 3 500 euro har man föreslagit för omedelbara kostnader - men vi uppmanar dem också att samarbeta på ett annat sätt med regeringen och de venezuelanska medborgarna .
Den här veckan talar vi också om en katastrof som inträffat i Europa och vi nämnde att de klimatologiska förändringarna kan ha haft något att göra med denna ökning av katastrofer som felaktigt brukar kallas naturkatastrofer , vilket redan har fastställts av många experter .
Vi tror att det är vi människor som bär skulden .
I Venezuelas fall - vi hade glädjen att vara där med anledning av konferensen mellan Europaparlamentet och det latinamerikanska parlamentet - är den brutala urbaniseringen och angreppen på miljön mycket märkbar och något som eventuellt kan förvärra sådana här situationer .
Herr talman , vi måste se till att infrastrukturen återuppbyggs .
De europeiska institutionerna , medlemsländerna , en del icke-statliga organisationer måste samarbeta med andra länder så att den här katastrofen , som orsakat irreversibla skador , kan mildras så gott det går .
Herr talman !
Jag är inte ute efter att vara övertydlig med tanke på tidigare anföranden , men jag kommer också från ett område , Baskien , där man känner stor solidaritet .
Venezuela har tagit emot emigranter från hela Spanien och då särskilt från Baskien och under de många och långa åren av diktatur fick vi ovärderlig moralisk och materiell hjälp .
Och eftersom " en olycka kommer sällan ensam " så har vi de senaste dagarna kunnat registrera såväl en jordbävning ( 6 grader på Richterskalan ) som en havsbävning .
Eftersom sorgen och solidariteten är delad vill jag centrera mitt anförande på en del frågor som ligger bortom det materiella biståndet på kort sikt och själva resolutionen .
Vi måste granska utvecklingsmodellen , inte bara Venezuelas utan också andra länders , och ta upp det som inte överensstämmer med bevarandet och respekten för miljön .
Bistånd måste avsättas även för detta ändamål och för den negativa inverkan en del industrisektorer står för i den ekologiska jämvikten , och inte bara i Venezuela .
Det är absolut nödvändigt att en konferens Europeiska unionen-Latinamerika hålls så att vi kan hejda tendensen av beroende och exporten av energiresurser samt den exploatering som i blindo sker av densamma .
Vi måste göra vad som står i vår makt för att förhindra katastrofer av det här slaget .
Frågor som dessa måste följaktligen uppmärksammas , men givetvis även dem som tas upp i resolutionen .
Avslutningsvis vill jag inte låta tillfället gå mig ur händerna utan att uppmärksamma angivelserna om kränkningar av de mänskliga rättigheterna i Venezuela under täckmanteln att hindra området från att plundras .
Vi får inte titta åt ett annat håll när det gäller det här heller .
Vår solidaritet med det venezuelanska folket får inte göra att vi blir mindre uppmärksamma på individer som president Chávez , en populistisk president som har visat prov på oroväckande intolerans och hot mot vissa sektorer , inklusive massmedia , även om det finns en del europeiska parlamentsledamöter som är beredda att " skratta åt hans lustigheter " .
I Venezuela bor mer än 300 000 av mina landsmän för att finna möjligheter till ett bättre liv .
Venezuela tog vänligt emot dem med öppna armar .
Det samma har skett med hundratusentals andra europeiska invandrare .
Jag kan för övrigt nämna att mer än 70 procent av de invandrade portugiserna i Venezuela kommer från min region , Madeira .
Denna stora närhet gjorde att vi följde katastrofen med djup sorg och sinnesrörelse .
Men den skapade också en stor solidaritetskänsla .
Det var därför mycket tacksamt att höra kommissionens meddelande om den humanitära hjälpen .
Emellertid har tragedins storlek visat hur otillräckligt denna hjälp är .
Sanningen är att Venezuela drabbats av den största naturkatastrofen i Latinamerika under 1900-talet .
Det är klarlagt att minst 15 000 människor har dött .
Hundratusentals har förlorat sina bostäder .
De uppskattade materiella skadorna uppgår till mellan 10 och 20 miljarder dollar .
Man har förlorat 230 000 arbetstillfällen .
Inför denna enorma och tragiska bild måste Europeiska unionen påtagligt öka sitt stöd till Venezuela .
I detta syfte har jag lagt fram detta resolutionsförslag i parlamentet .
Vi önskar att Europaparlamentet , de europeiska folkens representativa organ , reser dit för att visa sin sorg och solidaritet .
Vi vill också att parlamentet uppmanar kommissionen att stärka den humanitära hjälpen för att bidra till de oändliga behoven inom områden som sjukvård , vatten , offentlig hälsovård , livsmedelsförsörjningen etc .
Vi vill även föreslå kommissionen att utarbeta en handlingsplan på medellång sikt för återuppbyggnaden av infrastruktur och bostäder , eftersom återuppbyggnaden av katastrofområdet kan ta mer än sju år .
Denna plan måste prioritera och stimulera återupptagandet av den ekonomiska verksamheten genom ekonomisk stimulans , extra finansiering och specialiserat bistånd .
Vi vill också uppmana kommissionen att mobilisera så mycket som möjligt av nödvändiga medel för att kunna ta itu med det nämnda arbetet .
Vi vill inte bara nöja oss med goda intentioner .
Herr talman !
Detta är det minsta vi kan göra för den befolkning som har drabbats av översvämningarna .
Herr talman !
Jag menar att Europeiska unionen skulle begå ett stort misstag om vi undervärderade omfattningen av den tragedi som Venezuela upplevt och där , som vi har blivit påminda om , tusentals liv har gått förlorade .
Det är bra att vi uttrycker vår solidaritet , men det är viktigt och brådskande att vi går från ord till handling .
Gemenskapens svar bör vara ett vittomfattande projekt för återuppbyggnad och rehabilitering av landet och där olika aspekter beaktas : Att förstärka det humanitära stödet och det omedelbara stödet samt att inrätta rehabiliterings- och återuppbyggnadslinjer , som extra insatser .
När jag säger extrainsats så säger jag det därför att ministerrådet nästa måndag kommer att anta ett uttalande som baserar sig på ett avtal mellan Coreper-ambassadörerna vari man säger att bistånd skall ges efter förmåga .
Det är omöjligt att finansiellt prioritera detta med Mitch-resurserna .
Vad parlamentet ber om - och man ber om det som en av budgetmyndighetens två grenar - är att kommissionen lägger fram ett ambitiöst förslag som kan ge ett svar på den situation som uppstått .
Det vore intressant om kommissionen kunde granska såväl de möjligheter som en tillämpning av de kommersiella åtgärderna ger vid handen , inom det schema som förutses i det allmänna preferenssystemet , som en utvidgning och förlängning av Europeiska investeringsbankens krediter .
Som prov på vår solidaritet och vårt stöd borde Europeiska unionen också stödja en " internationell givarkonferens " .
Vi måste leva upp till de krav som denna lidande befolkning ställer på oss , de är Europeiska unionens vänner , liksom Venezuelas folk , och de förväntar sig detta av oss .
Herr talman !
Om man skulle projicera den skada som Venezuela har lidit på Tysklands territorium så vore det i stort sett det samma som om hela kustområdet hade förstörts och 200 000 människor hade omkommit .
Då förstår man vilka våldsamma dimensioner olyckan har fått för ett land som Venezuela .
Det är knappast makabert av mig att påstå att det bästa som för tillfället kan hända Venezuela är ett så högt oljepris som möjligt för att Venezuela skall kunna finansiera så mycket som möjligt av egen kraft .
Visst är det oangenämt för oss , eftersom det blir dyrt , men för Venezuela är det fördelaktigt .
I det avseendet har Venezuela trots all skada man har lidit det bättre förspänt än Mellanamerika hade efter orkanen Mitch .
Dock är detta en klen tröst i betraktande av den våldsamma ödeläggelsen .
Kraven på en internationell konferens med bidragsgivare under aktivt deltagande av kommissionen är därför av värde .
I övrigt väntar jag - liksom mina kolleger - på att kommissionen så snart som möjligt skall lägga fram en plan för hur man efter avstämmande med regeringen i Venezuela skall kunna hjälpa till .
Venezuelanerna litar på vår medkänsla .
Men de behöver givetvis även pengar , fantasi och medverkan vid återuppbyggnaden .
Tillåt mig att tillägga att globalisering faktiskt inte bara är handel utan även solidaritet .
Vid en så förhärjande katastrof är det naturligtvis även på sin plats att fråga efter orsakerna .
Jag är rädd att vi kommer att få sysselsätta oss allt mer med naturkatastrofer som människan är medskyldig till .
Visst , inför en naturlig klimatförändring står människan maktlös .
Men vid det här laget är växthusgaserna med i bilden .
Det är just där problemet ligger .
Tyvärr fullgör Europa inte sina förpliktelser från Kyoto .
Det är min förhoppning att denna katastrof - och tyvärr även andra - skall ge oss orsak att fundera över det här och att vidta åtgärder , så att de brådskande frågorna inte ständigt och jämt behöver handla om katastrofer , utan att vi kanske också kan diskutera vad vi i förebyggande syfte kan göra för att katastroferna inte skall bli så omfattande .
Om naturen nu kräver detta så bör människan åtminstone inte göra sig medskyldig .
( Applåder ) .
( FR ) Herr talman !
Kommissionen delar den oro som parlamentsledamöterna uttryckt för den katastrofala situationen i Venezuela och jag kommer att vidarebefordra era olika kommentarer till Nielsen .
Mot bakgrund av katastrofens omfattning reagerade kommissionen omedelbart genom att fatta beslut den 23 och 30 december 1999 , som redan nu genomförts , rörande beviljandet av en humanitär hjälp på 3,2 miljoner euro .
Med tanke på den omedelbara nödvändigheten att göra en utvärdering av behoven begav sig emellertid en expert från kontoret för humanitärt bistånd , ECHO till Venezuela redan den 22 december .
En ständig medarbetare från ECHO kommer att anlända till platsen inom de närmaste dagarna för att samordna den humanitära hjälpen och sköta genomförandet av programmen .
Med tanke på den höga risken för kolera- och spetälskeepidemier bland annat , som har bekräftats av hälsoministeriet i Venezuela , planerar kommissionen ett tredje beslut om 2 miljoner euro för att återställa ett dricksvattensystem och en epidemiologisk övervakning .
Jag delar Linkohrs åsikt beträffande tillfället att inför framtiden ha en allmän diskussion om katastrofer och vissa undersökningar går i den riktningen .
Utöver kommissionen svarade naturligtvis världssamfundet snabbt och generöst på regeringens vädjan .
Enligt FN : s Byrå för samordning av humanitär hjälp uppgår det sammanlagda beloppet för närvarande till omkring 24 miljoner dollar , varav nära 10 miljoner dollar från Europeiska unionen .
För att uppfylla parlamentets önskningar förbereder kommissionen emellertid också en expertresa för att bedöma situationen i Venezuela och identifiera speciella åtgärder .
Beroende på resultatet av expertutlåtandet kommer den att besluta om en uppbyggnadsplan på medellång sikt .
Kommissionen kommer att vara särskilt uppmärksam på frågor i samband med miljön när rehabiliteringsåtgärderna sätts in .
Vi är inte på det här stadiet i stånd att ange stödbeloppet , som kommer att bestämmas utifrån resultatet av expertutlåtandet och i samråd med andra givare .
Kommissionen skall ha ett nära samarbete med de övriga givarna för att uppmuntra till samordning av världssamfundets ansträngningar och fastställande av åtgärdsprioriteringar .
Det är således väsentligt att ett samordningssystem för den internationella hjälpen införs så snabbt som möjligt .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum kl .
17.30 .
( Sammanträdet avbröts fram till kl .
17.30 ) ( Sammanträdet avbröts återigen , från kl .
17.30 till kl .
18.00 . )
ORDFÖRANDESKAP : PROVAN vice talman Herr talman !
Jag vill att min protest förs in i protokollet , omröstningen skulle äga rum kl.17.30 och den har försenats utan någon som helst förklaring .
Det visar på bristande respekt mot kammaren och mot alla oss som var här till utsatt tid .
Detta kan bara rättfärdigas vid force majeur , som till exempel herr eller fru ordförandens hjärtinfarkt .
Om så inte är fallet anser jag detta visa på ett oförsvarligt förakt för oss parlamentsledamöter .
( Livliga applåder ) Herr Martínez !
Jag förstår er ståndpunkt fullständigt .
Allt jag kan säga er i detta skede är att detta kommer att hänskjutas till talmanskonferensen , som , själv , bad om fördröjningen .
Det är egentligen upp till plenum att fastställa föredragningslistan , men av en eller annan anledning beslutade talmanskonferensen , som fortfarande sitter i möte , att skjuta upp sammanträdet med ytterligare en halvtimme .
Jag lovar att se till att era anmärkningar vidarebefordras i de starkaste ordalag .
Jag hoppas att det tillfredsställer er alla .
Jag vill inte inleda en debatt om detta just nu .
Det är en sak som har skett .
Ju snabbare vi kommer igång med omröstningarna , desto bättre .
Låt mig försäkra er om att det är den sortens fråga som förtjänar en riktig diskussion och ett riktigt beslut av parlamentet självt snarare än ett enkelt ad hoc-beslut om att ändra föredragningslistan .
Under omröstningen om Tjetjenien Herr talman !
En synpunkt som gäller resolutionen om Tjetjenien .
Jag vill bara påpeka att det under punkt 4 i den tyska versionen talas om tjetjenska miliser , men i den engelska originaltexten talades det om fighter .
Fighter betyder emellertid stridskämpe .
Jag ber er alltså rätta till detta i alla språkliga versioner , därför att det är stor skillnad mellan fighter och miliser .
Under punkt 4 vill jag alltså be om granskning av de olika språkversionerna .
Ni har helt rätt , herr Posselt .
Texten kommer att anpassas i enlighet därmed .
Före omröstningen om Egypten Herr talman !
Jag ber om överseende , men det gäller återigen samma problem .
I den engelska originaltexten som låg till grund för förhandlingarna talas det om sectarian clashes eller något ditåt .
Hur som helst är det ordet " sectarian " det gäller .
I den tyska versionen heter det : " Strider mellan muslimska och koptiska sekter " .
Även detta är rena dumheterna , och jag ber er anpassa detta efter den engelska texten .
Återigen , vi kommer att se till att texten är korrekt översatt till tyska .
Efter omröstningen om Moluckerna ( Indonesien ) : Herr talman !
Den närvarande kommissionären sade att problemet med vapenembargot mot Indonesien troligen kommer att analyseras av rådets möte om allmänna frågor den 24 , vilket är på måndag .
Jag skulle alltså vilja be om särskild solidaritet från presidiet och stor omsorg att resolutionen vi har röstat igenom omedelbart sänds till rådet .
Och att sekretariatet ser till att handla mycket skyndsamt .
Jag tror att ministrarna läser tidningarna , men det är viktigt , eftersom det är andra gången Europaparlamentet uttalar sig för att förnya vapenembargot , att den resolution vi har röstat igenom omedelbart kommer till rådets kännedom .
Det skall ordnas .
Herr talman !
En ordningsfråga .
I morse lades två procedurmässiga förslag fram , ett av min kollega Hudghton och ett av mig själv .
Båda förslagen var förslag i vilka vi begärde en omröstning med namnupprop , för vi ansåg att det var angeläget .
Hittills finns i utskriften av omröstningarna med namnupprop endast namnlistan från den första , men inte - ännu - den andra , omröstningen om tillåtlighet .
Ledamöterna kommer nog ihåg att omröstning verkligen genomfördes med namnupprop och att den genomfördes med hjälp av maskinerna .
Kan vi garanteras att omröstningsrapporten kommer att finnas tillgänglig till i morgon bitti ?
Vi skall verkligen undersöka detta , herr MacCormick , och försöka se till att ni får den i tid att ta med den hem .
 
Den inre marknaden och rättsskydd för konsumenter Nästa punkt på föredragningslistan är debatt om den muntliga frågan ( B5-0039 / 99 ) av Palacio Vallelersundi för utskottet för rättsliga frågor och den inre marknaden till kommissionen om en balanserad strategi för den inre marknaden och konsumenternas rättsskydd .
Herr talman , herr kommissionär !
Eftersom vi har gått om tid vill jag ge ett exempel som kan vara lärorikt .
Det var en gång , innan Amsterdamfördragets ankomst , ett råd som debatterade en ändring av Bryssel- och Luganokonventionerna .
För dem som inte är förtrogna med teknikaliteterna så är det ett problem som berör domsrätten .
Med andra ord , inför vilken domare skall man beklaga sina sorger i en gränsöverskridande konflikt .
Rådet träffade en överenskommelse , enhälligt och inom ramen för det mellanstatliga samarbetet , det vill säga långt från gemenskapsandan men nära den internationella offentliga rätten .
Men plötsligt träder Amsterdamfördraget i kraft och i enlighet med artikel 65 var man tvungen att hantera ändringarna i Bryssel- och Luganokonventionerna som en gemenskapsfråga och de nya konventionerna omarbetas till en gemenskapsakt : en förordning .
Kommissionen tog då plats på scenen och mycket snabbt och för att skörda den första frukten av det nya Amsterdamfördraget bestämde man sig för att det räcker med att ändra rubrik för att omarbeta till en gemenskapsakt .
Där det står konvention skall det i stället stå förordning .
Därmed basta .
Kommissionen började således förbereda ett förslag till förordning om nämnda domsrätt , och detta utan att rådfråga någon , utan att rådfråga de olika generaldirektoraten .
I dag behandlar parlamentet betänkandet - fortfarande ett enkelt yttrande , eftersom parlamentet i den här frågan har begränsad behörighet - under ledning av Diana Wallis , som jag hoppas kommer att redogöra för det hela .
Av detta - och här slutar min historia - bör vi dra vissa slutsatser : För det första den bristande samordningen i rådet .
Rådet är inte rådet , det är rådet i betydelsen " rättvisa " .
Dessutom vill jag tillägga att det var en samling experter , professorer i internationell privaträtt , som förhandlade fram de internationella fördrag som , när allt kommer omkring , tar upp ämnet i fråga .
Man hade inte heller rådfrågat rådet ( inre marknaden ) och inte heller rådet ( allmänna frågor ) .
Även i kommissionen brast samordningen , vilket är viktigare för framtiden .
Förvisso höll kommissionen på att avgå och det var en svår period , men den bristande samordningen berodde faktiskt på att granskningen skedde efter det att förslaget till förordning hade offentliggjorts , varvid man gick emot alla elementära effektivitetskriterier och till och med respekten för medborgarna och kammaren , för att nämna något annat .
Det här exemplet visar också klart och tydligt vilken svår situation eller , herr talman , om ni så vill vilken stor utmaning vi står inför .
Kriterier för den inre marknaden , kriterier för den internationella privaträtten .
För att omarbeta en handling till gemenskapsakt är det verkligen bara fråga om att skriva förordning där det står konvention ?
Enligt utskottet för rättsliga frågor och inre marknaden så får det inte gå till på det viset och jag hoppas att parlamentet delar den uppfattningen .
För att omvandla en handling till gemenskapsakt måste man först och främst och framför allt göra en screaning av var och en av de normerande förslag som läggs fram i förhållande till den inre marknadens grundläggande principer .
Särskilt principen om ömsesidigt erkännande och principen om kontroll i ursprungslandet .
Att omvandla en handling till gemenskapsakt innebär faktiskt att vi visar respekt för den inre marknaden , vilket är mycket viktigt .
För att avsluta arbetet med den inre marknaden måste vi nämligen ta itu med de gränsområden som omger våra nuvarande lagar och eftersom de är förankrade i processrätten , och givetvis även i många delar av den internationella privaträtten , så finns här en klar definitionsbrist .
Om vi tappar bort de kriterier som håller den inre marknaden informerad tömmer vi indirekt meningen med denna och därmed styr vi in på en synnerligen farlig väg .
Det finns även en annan fara .
I den digitala revolution vi nu lever i finns en viss tendens att säga " vi är globala , den inre marknaden har blivit för liten , låt oss reglera världen , varför skall vi ha en inre marknad , låt oss hoppa över den " .
Nåväl , kom ihåg att den europeiska integrationen byggdes på den inre marknaden och att vi dessutom genom ett fördrag är förbundna att respektera de principer som stöttar och gestaltar denna verklighet .
Var finns då konsumenterna , frågar ni mig .
I det exempel jag gav så är det faktiskt så att man försöker skydda dem genom att ge dem en möjlighet att gå till domaren i grannhuset och be honom skipa rättvisa , gå till en domare där man har sin hemvist .
Är detta att skydda dem ?
Nej , det är det inte .
Ett bevis på detta är att konsumenterna inte processar när de köpt en liten sak , när de köper en liten sak i närbutiken .
Varför ?
Därför att det är mycket dyrt och tar väldigt lång tid .
Vill vi skydda konsumenterna måste vi vidta åtgärder .
Till exempel de två som kommissionen presenterat , small claims procedure eller ett utomrättsligt förfarande vid konsumentkonflikter .
Detta skyddar konsumenterna : Snabba , billiga och effektiva förfaranden .
Dessutom , herr talman , så skyddar vi konsumenterna genom att behandla dem som vuxna och inte tro att de är människor som inte klarar av att välja .
En av Europas största utmaningar i dagens digitala revolution är enligt min mening att ändra kulturen och rådande principer i konsumentskyddet .
Konsumenterna måste skyddas , de måste skyddas i verkligheten , inte bara formellt , och en riskfaktor måste tas med i beräkningen , en för konsumenterna beräknad risk så att de fullt medvetna kan göra sitt val .
Herr talman , snart slutar jag .
Europa måste försvara sina värden , men Europa står också inför en annan stor utmaning , jämvikten mellan den offentliga lagstiftningen och self regulation .
För att skydda konsumenterna måste vi ha en solid och skyddande ram för den offentliga lagstiftningen , men vi behöver också ett utrymme så att vi från det civila samhällets sida kan inrätta system som bättre passar in i den tid vi lever än vad de offentliga institutionerna kan göra .
Vid toppmötet häromdagen i Madrid sade någon till mig : " Fru Palacio , med Internet är ett år som två månader .
Ett direktiv som ni tar fyra år på er att fastställa är en väldigt lång tid " .
Låt oss skynda på , låt oss bevara våra värderingar men vi måste förstå att den inre marknaden är en prioritet . .
( NL ) Herr talman !
Jag skulle gärna vilja börja med att tacka ledamoten , Palacio , som ger mig möjlighet att gå in på ett ämne som är utomordentligt viktigt och även utomordentligt komplext .
Jag skulle vilja säga följande om det .
Liksom Palacio fäster kommissionen , med tanke på åstadkommandet av ett område utan inre gränser , som avses i artikel 2 i Fördraget om Europeiska unionen , stor vikt vid principen att företag skall kunna erbjuda sina varor och tjänster i hela unionen utan att den berörda medlemsstaten skall kunna sätta upp diskriminerande och orättvisa hinder .
Sådana hinder kan nämligen leda till en splittring av den inre marknaden genom att företag måste anpassa sina varor och tjänster till föreskrifterna i alla de EU-länder som de är verksamma i .
Det är vår utgångspunkt .
Det är en utgångspunkt som Palacio delar .
Hon sade för övrigt alldeles nyss att Europeiska unionen grundar sig på den inre marknaden .
Det håller kommissionen fullständigt med Palacio om .
Villkoret för ett fullständigt godkännande av principen om ömsesidigt erkännande är dock att alla medlemsstater har en lämplig och jämförbar nivå av konsumentskydd .
I det förslag till direktiv angående vissa juridiska aspekter av den elektroniska handeln som ledamoten nämnde anges tydligt att begreppet " inre marknad " i artikel 3 inte omfattar förpliktelser i konsumentavtal .
Som Palacio vet så regleras förpliktelser i konsumentavtal genom Romkonvention I och det är alltså fristående från det direktiv om elektronisk handel som rådet nådde politisk enighet om den 7 december förra året .
När det gäller de nyligen framlagda initiativen från kommissionen inom ramen för den nya avdelningen IV i Fördraget om upprättandet av Europeiska gemenskapen så antar jag att Palacio framför allt , och det sade hon egentligen också alldeles nyss , avser det förslag till förordning som kommissionen godkände i juli 1999 , på grundval av verksamheterna i en ad hoc-grupp i rådet och efter det politiska godkännandet från de femton medlemsstaterna , och vars syfte är att i gemenskapsrätten införliva Brysselkonventionen från 1968 angående domstols behörighet och verkställighet av domar inom det privat- och handelsrättsliga området .
Palacio tog upp det som hastigast och hon kritiserade det sätt på vilket kommissionens föreslagna förordning kommit till .
Hon sade också att det inte förekommit mycket samråd , inte bara mellan kommissionen och parlamentet utan till och med inbördes mellan de olika råden .
Kommissionen föreslog ändringarna och det ursprungliga avtalet från 1968 för att anpassa det redan gamla avtalet till moderna handelsmetoder och framför allt till elektronisk handel .
Nu verkar ledamoten anse att utgångspunkterna för det här förslaget till förordning , vilket alltså skall införliva Brysselkonventionen i gemenskapsrätten , skulle kunna vara i strid mot principen om ursprungslandet .
Det skulle emellertid , om hon hade rätt , innebära att även domstols behörighet skulle omfattas av den principen och det är inte fallet .
För övrigt anges det i artikel 1 i det nämnda förslaget till direktiv om elektronisk handel , såsom det fastställdes i en politisk överenskommelse i december , att det förslaget inte gäller för frågan om domstols behörighet .
Som Palacio vet så omfattas frågan om domstols behörighet av Brysselkonventionen .
Situationen i dag är alltså den att det finns tre parallella akter .
Det finns ett föreslag till direktiv om elektronisk handel .
Vi har Romkonventionen som jag nyss hänvisade till och vi har Brysselkonventionen .
Det är tre akter som just nu existerar oberoende av varandra .
Kommissionen skall se till , herr talman , att det på lämpligt sätt tas hänsyn till de invändningar som främst yttrades vid utfrågningen den 4 och 5 november , angående eventuella effekter av det här förslaget till förordning för den inre marknaden samt även till de förklaringar till förmån för förslaget som mottagits .
Kommissionen analyserar just nu de mångfaldiga och detaljerade ståndpunkter som den mottagit och skall i sinom tid tillkännage eventuella förslag .
I varje fall verkar det dock vara önskvärt , särskilt i ljuset av den kritik som Palacio fört fram , att kommissionen , innan den tar något initiativ , först känner till den ståndpunkt som Europaparlamentet i februari i år skall anta angående förslaget .
Det verkar också vara nödvändigt att lämpliga , kompletterande lösningar hittas för att tillmötesgå de invändningar som lades fram av konsumentföreträdare vid utfrågningen .
Därför måste förhandlingar snabbt inledas med alla berörda parter för att komma fram till alternativ , vilket även Palacio bett om , till de ofta långdragna , dyra och invecklade rättsprocesserna för att snabbt och mindre dyrt för konsumenten avgöra tvister som uppstått på grund av elektronisk handel .
Herr talman !
Låt mig först av allt tala om hur mycket jag välkomnar det som Bolkestein just har sagt om att kommissionen skall genomföra en mycket ingående granskning av de komplexa och överlappande lagstiftningsdelar som kommer att påverka den nya värld som vi lever i - den elektroniska handelns nya värld .
Jag hade turen att kunna närvara på delar av utfrågningarna den 4 och 5 november , och antalet inblandade människor och kvaliteten på bidragen visar hur allvarligt folk tog frågan .
Det är en återspegling av den oro som fanns över det ursprungliga synsättet .
Min kollega Wallis , som utarbetar vårt betänkande , kommer att tala om en stund , och jag vill inte föregripa eller stjäla det som han skall säga .
Vi kommer att diskutera det senare , och jag vet , herr kommissionär , att ni redan har sett några av delarna i det .
Den punkt som jag vill ta upp skall jag inte ta upp med en jurists perspektiv , eftersom jag har privilegiet att vara en av de få i utskottet för rättsliga frågor och den inre marknaden , under Palacios ordförandeskap , som inte är jurister .
Jag skulle vilja anlägga ett perspektiv på frågorna ur både handelns och konsumenternas synvinkel .
Nyckelordet i denna fråga som vi ställer till er , herr kommissionär , är balans .
Om vi ser oss runt i världen , håller ankomsten av elektronisk handel eller elektronisk kommunikation påtagligt på att ändra balansen på marknadsplatsen .
Balansen rör sig i en riktning som kraftigt gynnar konsumenterna .
Vi håller alla på att bli informerade konsumenter , eftersom den nya kommunikationstekniken ger oss enorma möjligheter att handla globalt , jämföra priser och fatta våra beslut på grundval av stora mängder lättillgänglig information .
De av er som inte har prövat på det , borde verkligen göra det , eftersom den elektroniska handeln , tack vare denna kombination av datorkraft och information , gör det möjligt för människor att jämföra erbjudanden och handla på ett sätt som de aldrig tidigare har gjort .
Jag skall ge er ett enkelt exempel .
Det är ett exempel som är av betydelse för vårt lagstiftningsarbete i hela den offentliga sektorn .
Telekommunikationsverket i Storbritannien har en webbsida som konsumenterna kan besöka för att jämföra detaljerna i de olika telekommunikationsbolagens erbjudanden .
Man skriver in detaljer om sitt telefonanvändande och jämför därefter de olika erbjudandena - det är den sortens möjligheter som inom kort kommer att vara tillgänglig för oss .
Denna nya generation av informerade konsumenter kommer inte att bekymra sig om argument som vi kan ha som lagstiftare om rättsprinciper och lagars tillämplighet , eftersom , vilket Palacio påpekade , rättsskydd inte är det som mest upptar tankarna hos människor som handlar , på Internet eller någon annanstans .
Innan ett beslut fattas om ett köp , kommer kunderna att vilja vara säkra på att den organisation som de har att göra med erbjuder bra villkor och garantier samt tillgång till tvistlösning .
Om det rör sig om ett relativt okänt märke - och vi bör uppmana små företag att använda den elektroniska handeln för att nå ut till konsumenterna - kan dessa konsumenter mycket väl vilja ha den trygghet som någon slags godkänt märke , ett e-handlarmärke , erbjuder , som till exempel det som den brittiska konsumentföreningen verkar för med stor framgång .
Vi måste berömma dem för det .
Det är den sortens initiativ vi måste uppmuntra runt om i Europeiska unionen .
Det är någonting som jag skulle vilja be kommissionären att ta upp som en del av denna serie frågor som hör samman med konsumentlagstiftning .
Människor kommer att vilja ha att göra med organisationer som hanterar problem och klagomål med samma hastighet och effektivitet som de gör sitt köp på Internet .
De kommer att vilja ha en enkel och effektiv tillgång till tvistlösning och tillgång till någon som kan hjälpa dem med deras problem En sak är säker om den elektroniska handeln , och det är att den verkligen utvecklas mycket snabbt .
Nya former av produkter och tjänster kommer ut på marknaden mycket snabbare än någonsin tidigare , och vårt jobb som lagstiftare i detta parlament är att uppmuntra denna dynamiska kraft , inte att dämpa den .
Vi vill uppmuntra konsumenterna att använda elektronisk information som underlag för sina köpbeslut och uppmuntra företag av alla storlekar , särskilt de små företagen , att delta i den elektroniska handeln .
Det kommer helt klart att göra det nödvändigt för oss att ompröva vårt regelverk .
Herr talman , ärade kommissionär !
Vi fortsätter i dag debatten om en balanserad strategi för den inre marknaden och rättsskydd för konsumenter på grundval av en muntlig fråga som framför allt behandlar motsättningen mellan principen om ursprungsland på den inre marknaden och principen om bestämmelseland i konsumentskyddet .
För muntliga frågor är dylika avkortningar oundvikliga .
Jag anser dock - vilket debatten hittills också har visat - att diskussionen om dessa bägge principer egentligen inte leder oss vidare här , särskilt inte när det handlar om att finna en lämplig rättslig ram för trafiken med elektronisk handel .
Det är med rätta man befarar - det medges - att konsumenternas möjlighet att i hemlandet väcka åtal enligt inhemsk lag kan ha en hämmande eller rentav avskräckande inverkan på etableringen av den elektroniska handeln .
Samtidigt vet vi emellertid också att möjligheten att väcka åtal på nationell bas ofta bara är en teoretisk möjlighet som inte utnyttjas .
Än mindre kan vi begära att konsumenterna skall behöva väcka åtal i leverantörens ursprungsland med följden att leverantörerna slår sig ned i de medlemsländer som har sämst villkor för konsumentskydd och där det svagaste rättsskyddet för konsumenterna anammas .
Det nödvändiga förtroendet från konsumenterna , vilket den elektroniska handeln ju också behöver för att utvecklas , blir säkerligen inte starkare av detta .
Därför tror jag egentligen inte att vi är hjälpta av vare sig den nya artikeln 15 i förordningen som sådan eller av dess begränsning till offline-affärer .
Vad vi saknar är system för biläggande av tvist utom rätta och metoder för att snabbt klara upp alla berömda small claims .
Därför välkomnar jag verkligen de åtgärder som kommissionen har föreslagit i sitt meddelande om framtida strategi , i synnerhet bidraget med initiativ till metoder om biläggande av tvist utom rätta , vilka tillämpas online , och till en ny grönbok om konsumenternas möjligheter när det gäller lag och rättsliga medel .
Dock anser jag att det också borde vara möjligt att tillsammans med de europeiska bankerna och kreditkortsleverantörerna utveckla en säker elektronisk penningtrafik liksom gireringssystem som möjliggör elektroniska steg för steg-affärer .
Även ett förstärkt samarbete mellan konsumentskyddsorganisationerna och gränsöverskridande befogenheter för dessa konsumentskyddsorganisationer skulle i slutändan vara oss mer behjälpliga i vardagen än en teoretisk tvist mellan bestämmelselands- och ursprungslandsprincipen .
När nu kommissionens preliminära förslag till ny förordning har kritiserats här vill jag med eftertryck påpeka att jag håller kommissionens tillvägagångssätt för korrekt .
Redan nu regleras i artikel 13 i konventionen hur domstols behörighet för konsumenter ser ut , redan nu tenderar den huvudsakliga åsikten bland jurister vara att detta gäller även för handel online .
Kommissionen ändrar här alltså ingenting i det aktuella rättsliga läget .
Och enligt artikel 95.3 , måste kommissionen som bekant utgå från en hög konsumentskyddsnivå .
Därför anser jag att kommissionen har agerat riktigt med sitt förslag .
Vi i den socialistiska gruppen stöder även förslagen från Wallis i utskottet för rättsliga frågor och den inre marknaden , som har föreslagit ett par ändringar i förslaget till förordning , men som även insisterar på att vi skall komplettera det aktuella systemet för att få fram nya metoder .
Jag vill avslutningsvis tala för min grupp och säga att det för oss är tänkbart att övergå till principen om ursprungsland endast om detta åtföljs av kravet på stärkt rättsskydd för konsumenten via nya metoder som ger möjlighet till rättsligt skydd .
Herr talman !
Med denna fråga uppmärksammas den spänning som finns mellan företagens och konsumenternas intressen inom ramen för den inre marknaden - en spänning , måste jag säga , som jag har blivit allt för bekant med som föredragande för Brysselkonventionen .
Idén om samordning har nämnts .
Jag vill fästa uppmärksamhet på en modell , eller kanske ett modeord , om ni så önskar , som för närvarande används mycket i Förenade kungariket angående styrelseformer .
Vi talar om sammankopplat tänkande eller sammankopplad förvaltning .
Det rör sig , med andra ord , om att överbrygga klyftor mellan departementen .
Detta är också ett mognadstecken , som när vi i skolan gradvis övergår från att texta till att använda skrivstil ; det vill säga vi kopplar samman bokstäverna .
Debatten om jurisdiktion och elektronisk handel har belyst denna konflikt mellan konsumenter och webbförsäljare .
Kan en konsument väcka åtal i sin egen domstol , om han är berättigad till det ?
Kommer detta att vara dödsstöten för den elektroniska handeln ?
Jag föreslår ett åtgärdspaket , i vilket frågan om rättsskydd , som vi hörde mycket om i Tammerfors , är central .
Om det inre marknaden skall fungera bra - om den fullt ut och med förtroende skall utnyttjas av både små företag och konsumenter - måste det finnas ett rättsskydd i civilrättsliga ärenden .
Det måste finnas förfaranden för små tvister och alternativa metoder för tvistlösning .
Det är absolut nödvändigt för den inre marknaden .
Men vår kommissionär kommer naturligtvis att säga att detta kanske ligger mer på hans kollega Vitorinos , och kanske också Byrnes , område .
Detta har frustrerat mig .
Byrne och Vitorino har talat om att upprätta system för lösning av små tvister i Europa .
Vi måste sammanställa dessa uttalanden till en helhet .
Kommissionen måste börja tänka på ett sammankopplat sätt - som en sammankopplad förvaltning .
Vi har ett en-chans-på-generationen-tillfälle att underlätta den elektroniska handelns tillväxt .
Angående den andra frågan , vi tycks i ökande utsträckning se harmonisering som ett sätt att lösa vissa av dessa problem - att lösa de spänningar som har uppstått .
Men det är ofta denna harmoniseringsprocess , som i alltför hög grad kan vara beroende av lagstiftning , som kan vara stel och inflexibel och som sedan själv blir en barriär mot den inre marknaden .
Det har hörts sådana påståenden om dataskyddsdirektivet , som är en viktig del av konsumentskyddslagstiftningen , men det verkar som om direktivet i vissa medlemsstater har tillämpats i överdriven utsträckning , vilket har lett till en potentiell barriär inom den inre marknaden .
Den elektroniska handeln är i mångt och mycket en global marknad .
De lösningar som vi antar måste tillåta våra medborgare och företag att delta på denna större marknad .
I Amerika - som inte nödvändigtvis måste vara vår förebild - har man valt en kombination av självreglering och mjuk lag uppbackad av lagstiftning .
Vi bör vara beredda på att undersöka denna slags blandning av lösningar .
En har redan nämnts .
En möjlig lösning kan ligga i kreditkortsindustrins händer .
Men för att kunna använda dessa lösningar , måste vi agera , och kommissionen måste agera gemensamt på ett sammankopplat sätt .
Herr talman !
Jag skulle vilja tacka Palacio och Bolkestein för att de har inlett denna diskussion med sedvanlig klarhet och hövlighet .
Det är anmärkningsvärt - och även om det kanske är banalt att säga det , kan jag inte låta bli - vilken enorm förändring den elektroniska handelns utveckling kommer att innebära för våra liv under de kommande årtiondena och under detta århundrade .
Vad beträffar mig själv , julhandlade jag på webben för första gången nu i julas , delvis på grund av de nya omständigheterna i mitt liv och min sämre tillgång för närvarande till köpstråken i Edinburgh .
Jag sände faktiskt blommor via elektronisk handel till min dotter på hennes bröllop nyligen i Texas , och som ni säkerligen förstår , herr talman , var det trevligt för en skotte att få blommorna dit utan någon biljettkostnad !
Vi rör oss in i en ny värld .
Men det finns , vilket har påpekats , utomordentligt svåra problem på detta område .
Om man ser bortanför det egna landet , kommer små företag att ha svårt att ta sig in på marknaden .
Berger tog upp en del av detta problem , men är det inte viktigt att komma ihåg att människor som ger sig in i affärer måste veta vad de behöver gardera sig mot , och lokal rådgivning om detta kommer att bli bättre .
Det gör det viktigt att hemlandsprincipen gäller .
Men sedan finns även det motsatta problemet .
Vi kan få se uppskörtningar på distans av företag i andra länder som vet att det inte är särskilt stor risk att de behöver möta arga fru Smith som har fått en oduglig vara med posten .
Hur tar man itu med det ?
Det har redan sagts två gånger - och det är en viktigt uppslag - att det borde finnas sätt att använda kreditkortsföretagen som en riskspridningsmekanism , under förutsättning att de är villiga att delta .
Konsumenterna kan ha rättigheter gentemot kreditkortsföretaget i sitt eget land , och kreditkortsföretaget kan ha rättigheter gentemot producenten eller säljaren i det landet .
På så sätt skulle alla de som agerar på marknaden delta till en liten del i riskerna över hela marknaden .
Kommissionen bör undersöka detta .
På lång sikt måste vi emellertid röra oss mot en harmonisering av lagarna för civilrättsliga och kommersiella ärenden i hela unionen .
Vi i Förenade kungariket hade , som ni känner till , herr talman , en mycket framgångsrik inre marknad under 300 år , med två rättssystem som växte ihop spontant , inte genom tvång .
Vi måste i det långa loppet sträva mot den typen av utveckling i Europa .
Vi borde ha europeiska riktlinjer som de amerikanska riktlinjerna och låta våra lagar utvecklas .
Herr talman !
Jag företräder en ståndpunkt som jag delar med Nobilia , tillsammans med vilken jag ingår i en speciell grupp inom UEN-gruppen .
Vi anser att det problem som tagits upp av Palacio förmodligen är ett av de viktigaste problem som den inre marknaden står inför .
Lagstiftningen på detta område är bristfällig och senfärdig och i stället för att erbjuda konsumenterna en grundsäkerhet och ett enhetligt rättsligt skydd , så lämnar den stora marginaler för ogrundat godtycke och oklarheter .
Detta gäller utan tvekan det område frågeställaren angav som ett exempel - den elektroniska handeln - och i samband därmed försäljningsmetoderna , köparens rättigheter , möjligheterna att få rättelse och också de olika skattesatser som tillämpas på själva försäljningen .
Men problemet kommer även att beröra oräkneliga andra områden : till exempel elektroniska komponenter , där produktionen kan ske i flera olika länder , även utanför gemenskapen , lagring och / eller anbringandet av varumärket kan ske i en medlemsstat och slutmonteringen i en annan .
Problemet gäller inte så mycket de olika komponenterna pålitlighet och om man respekterar lagstiftningen i import- eller tillverkningslandet , utan snarare hur de i sin helhet ger en ökad flexibilitet .
Detta är synpunkter som får ett kraftfullt stöd inom Europeiska unionen , framför allt om de länder där produktens slutlige konsument är bosatt , i avsikt att uppnå en bättre konkurrenskraft för de ekonomiska aktörer som verkar inom landet , har inrättat ett system med ursprungsbeteckningar som utgår från klart angivna egenskaper som bestämts tidigare och som går utöver det som bestämts av unionen .
Detta är något som framför allt förekommer inom livsmedelsproduktionen , där problemet , som framför allt rör ursprungslandet , som en följd av de undantag som medlemsstaterna beviljats i detta avseende , i första hand uppkommer i samband med den information som skall lämnas på etiketten till den produkt som är avsedd att gå till den slutlige konsumenten .
Det är uppenbart att en sådan situation inte bara skapar obeslutsamhet och osäkerhet utan samtidigt ändrar konkurrensförhållandena till nackdel för de små och medelstora företagen , inte när det gäller respekten för den ena eller andra nationella lagstiftningen , utan när det gäller de försämrade möjligheter de får på grund av brister i gemenskapslagstiftningen .
Det är också uppenbart att om dessa nackdelar för de små och medelstora företagen får fortsätta kan man frukta återverkningar på sysselsättningen , som man inte kan undvika vare sig genom att förenkla de administrativa rutinerna eller genom att minska företagsbeskattningen , eller genom att engagera arbetsmarknadens parter och deras resurser .
Detta innebär att man vid sidan om arbetet med att utarbeta särskilda förordningar för de produkter och de speciella förhållanden som angetts ovan , också måste förstärka den gemensamma vision och lagstiftningsfilosofi som krävs för att skapa ett riktigt regelsystem för den inre marknaden , ett regelverk som kan bli en effektiv referenspunkt och skapa trygghet för medlemsstaterna och för alla ekonomiska aktörer .
Avslutningsvis anser vi att det vid sidan om den kontroll av fragmenteringsgraden som kommissionen genomfört - ett verkligen berömvärt arbete när det gäller tillnärmningen av den nationella lagstiftningen - så måste man även göra alla ansträngningar för en korrektare tillämpning och en snabbare överföring av det mandat som rådet i Wien gav , och som sedan dess understrukits just när det gäller den inre marknaden , för att förbättra den europeiska ramlagstiftningen och konkurrenskraften , något som mycket väl kan få åtföljas av undanröjda handelshinder och en effektivare administration .
Herr talman !
Den muntliga frågan från utskottet för rättsliga frågor och den inre marknaden med avseende på eventuella handelshinder som kan uppstå genom konsumentlagstiftning innehåller redan en lösning på dem : ytterligare harmonisering .
Men behövs det verkligen ?
Genom den inre marknaden har det blivit lättare för producenter och konsumenter att ta steget över gränsen .
För sådana gränsöverskridande transaktioner behövs det en lämplig lagstiftning .
Därför behövs det en minsta harmonisering av lagstiftningen .
En hög nivå av konsumentskydd betyder inte att allt måste regleras europeiskt genom maximimal harmonisering .
Tvärtom , vi måste söka efter den bästa lösningen för konsumenten , i det här fallet en tillförlitlig referensram .
Det kommer ofta att vara en nationell ram .
Vid elektronisk handel kan ursprungsland väljas ganska godtyckligt .
Det är inte bra för konsumenternas förtroende .
Därför måste konsumenten få möjlighet att välja det egna landets lagar .
Att det skulle ge oönskade handelshinder tycker jag inte verkar rätt .
Konsumentskydd skapar en nödvändig , politiskt önskvärd förutsättning för handeln , till skydd för den svagare parten .
Kommissionens handlingssätt leder i varje fall inte till en ändlös dragkamp om önskvärd harmoniseringsnivå .
Det kräver inte heller någon ny lagstiftning på gemenskaps- eller nationell nivå och subsidiaritetsprincipen respekteras .
Det finns inget obalanserat i kommissionens strategi .
Möjligen i det utskottets för rättsliga frågor , som ständigt hamrar vidare på gemenskapsstödet med argument som jag tycker är ovidkommande .
Herr talman !
En topprioritet för Europeiska kommissionen och även en topprioritet för den europeiska industrin och handeln är e-commerce , elektronisk handel .
Vi får inte glömma bort att även konsumenten har stor nytta av att på ett bra sätt kunna använda sig av e-commerce .
Vad kan vi nu konstatera ?
Det pågår en häftig diskussion mellan näringsliv och konsumenter om vilken rätt som skall tillämpas vid gränsöverskridande handel , vilket i allt högre grad omfattar den elektroniska handeln .
De som säljer varor och tjänster är för ursprungslandsprincipen , enligt vilken den lag som gäller i det land den som erbjuder tjänsterna och varorna är etablerad i skall tillämpas .
Det kan jag mycket väl förstå .
Herr talman !
Ett exempel .
En portugis köper en dator från Finland via Internet .
Finländarna har för övrigt ett mycket bra konsumentskydd .
Då gäller alltså ursprungslandsprincipen enligt finländsk rätt .
Den dyra datorn kommer dock inte fram fast du redan har betalt med ditt kreditkort .
Skulle den här portugisen vilja inleda en rättsprocess i Finland ?
Det tror jag inte .
Det skulle innebära att du också måste skaffa juridisk rådgivning i Finland eller om det finländska rättssystemet .
Det är dock inte allt , herr Bolkestein , det finns mer .
Mer än det som ni tagit upp .
Den europeiska konsumenten skyddas nämligen genom fler regler än endast de regler som gäller e-commerce eller de förordningar som ni nyss nämnde .
Det finns nämligen också ett direktiv om " distansförsäljning " .
Det kommer ett direktiv om " finansiella tjänster " .
Det finns också ett direktiv om privacy .
Där finns alla konsumentens minimivillkor och ibland även maximivillkor .
De föreslagna reglerna för e-commerce innebär att ytterligare ett antal extra åtgärder tillfogas .
Det finns två olika kommissionsförslag angående den här punkten .
Åtminstone angående rättsskyddet , nämligen vem kan man vända sig till ?
Å ena sidan alltså e-commerce som grundar sig på ursprungslandsprincipen och å andra sidan förslaget till den nya anpassade förordningen från Bryssel .
Jag håller dock med Bolkestein om att även om båda förslagen bokstavligen helst borde kombineras så är den bakomliggande tankegången dock motstridig .
Det leder alltså till förvirring och därför hindras det rättsliga skyddet vid e-commerce från att komma i gång på riktigt .
Herr talman !
Jag tycker att vi som Europaparlament borde ta ansvaret för att skapa ett bra konsumentskydd .
Konsumenten har nytta av ett genomblickbart och konsekvent system för rättsligt skydd .
Utan konsumenternas förtroende kan e-commerce nämligen inte riktigt gå sin egen väg och utvecklas fullt ut .
Därför måste vi , tycker jag , i högre grad än vi tidigare gjort , tänka : vilka är nu de alternativa möjligheterna för att ge konsumenten ett rättsligt skydd , även när något går fel ?
Då tror jag , och därför vänder jag mig även till kommissionär Bolkestein , att vi mycket hellre borde undersöka de alternativa systemen för avgörande av tvistemål .
I Nederländerna har vi , som ni vet , ett mycket välbalanserat system för alternativa avgöranden av tvistemål .
Det systemet är för övrigt mycket väl lämpat för gränsöverskridande ärenden varvid de instiftade tvistemålskommittéerna gör det möjligt för personer från utlandet att komma till Haag och protester vid de här kommittéerna och att även rättvisa skipas där .
Herr talman !
En av lösningarna är : börja leta efter en annan kurs att slå in på .
Herr talman , mina damer och herrar , kära kolleger !
Låt mig först tacka Palacio Vallelersundi för initiativet till en muntlig fråga .
Vad handlar detta om ?
Som slagord låter sig problemställningen omskrivas som följer : Konsumentskydd och elektronisk affärsverksamhet i hetluften .
Eller annorlunda uttryckt : Hur kan konsumenterna i Europeiska unionen skyddas effektivt utan att detta hindrar utvecklingen av e-commerce ?
Diskussionen koncentreras för tillfället till frågan om enligt vilken princip domstols behörighet och i förlängningen den tillämpliga lagen skall fastställas vid gränsöverskridande tvister inom den elektroniska affärsverksamheten .
Måste inte en konsument i ett tvistemål driva igenom sina rättigheter i det land där leverantören av varor eller tjänster har sitt säte , eller i det land där han bor ?
Vilken lag är det som skall tillämpas ?
Jag skall inte ta upp argumenten för och emot i dessa frågor igen .
Dessa aspekter är kända nog .
Kommissionen genomförde en hearing angående detta i november .
Jag vill i dag bara rikta uppmärksamheten på att diskussionen konsumentskydd å ena sidan och e-commerce å andra sidan enligt min mening förs för snävt , för korthugget .
Den står också i strid med strategin så som kommissionen själv har formulerat den i sitt meddelande om strategi för den inre marknaden .
I meddelandet från kommissionen förklarar man uttryckligen att balanserade lösningar skall finnas ifall konsumenternas och näringslivets intressen går isär .
Därvid skall utvecklingen av elektronisk handel i Europeiska unionen ges en realistisk chans .
Men en balanserad lösning står att finna i spänningsfältet mellan konsumentskydd och e-commerce business endast om diskussionen inte begränsas till frågan om domstols behörighet och tillämplig lag , utan i stället förs på bred bas .
Målet med överläggningarna om ett effektivt konsumentskydd måste ju vara att konsumenten på ett snabbt , kostnadseffektivt och obyråkratiskt vis skall kunna få ut sin rätt .
Förhåller det sig verkligen så när konsumenten på hemorten kan väcka åtal på grundval av lagen i det egna landet ?
I och med en dom i hemlandet ger man konsumenten i princip bara stenar för bröd , eftersom han måste verkställa eller fullborda sin dom i annat medlemsland .
Detta blir ofta utdraget , mödosamt och kostnadsintensivt .
För ett effektivt konsumentskydd måste det till en utvärdering av alternativ till kostsamma och tröga domstolsförfaranden , vilken domstol och vilken lag det än må gälla .
Biläggande av tvist utom rätta , i förekommande fall knutet till fortsatt standardisering , är enligt min mening det magiska ordet .
Generaldirektoratet har redan ingående behandlat frågan om utomprocessuell förlikning i samband med gränsöverskridande ekonomiska tjänster .
I oktober förra året genomfördes en hearing på detta tema .
Jag vill föreslå att insikterna och idéerna i kommissionens diskussionsunderlag , vilket låg till grund för hearingen , samt det meddelande om resultaten från hearingen som väntas kring halvårsskiftet utvärderas i detalj även för den elektroniska handeln .
Denna början till riktlinjer för e-commerce är enligt min åsikt politiskt sett mer fördelaktig och får därför inte omintetgöras av regleringen i Bryssel / Lugano-konventionen och i Rom II .
Därför föreslår jag inför det fortsatta arbetet antingen att ändringen från Bryssel / Lugano skjuts upp tills alla öppna lagfrågor på detta område har retts ut , eller också att status quo i intresseutjämningen mellan leverantör och konsument bibehålls när man ändrar Bryssel / Lugano . .
( NL ) Herr talman !
Jag skulle gärna i korthet gå in på några av de viktiga punkter som parlamentsledamöterna tagit upp .
Jag vill börja med ett uttryck som Harbour använde och jag skulle också vilja ta tillfället i akt att tacka herr Harbour för det stora intresse han visade vid frågestunden den 4 och 5 november .
Kommissionen uppskattar det alltid väldigt mycket när parlamentsledamöter deltar vid en frågestund och andra verksamheter , och jag skulle gärna vilja understryka det här , herr talman .
Harbour talade i alla fall om jämvikt och det är naturligtvis det som kommissionen eftersträvar .
Ni skall förstå , herr talman , att jag inte bara talar för min egen del och för mitt generaldirektorat utan även för hela kommissionen .
I kommissionen sitter bland andra min kollega Byrne , som handhar konsumenternas intressen , och i mina svar vid den här debatten måste jag naturligtvis också ta hänsyn till Byrnes ståndpunkter så att vi , som Wallis kallade det , uppvisar en joined up-administration .
Den jämvikten eftersträvar vi och det är en jämvikt mellan å ena sidan producentens intressen och å andra sidan konsumentens intressen .
Det är välkänt och även argumenten är naturligtvis tydliga .
Den jämvikten eftersträvar vi .
Jag tror att vi lyckats uppnå den jämvikten i direktivet avseende elektronisk handel .
Principen i direktivet är att ursprungslandet spelar en avgörande roll när det uppstår tvister i samband med elektronisk handel .
Det är en avvikelse från den allmänna ordningen , så skulle jag kunna formulera det .
Den avvikelsen är dock mycket noga angiven .
Det måste handla om vissa ändamål och inga andra .
Det måste vara en avvikelse som är nödvändig .
Landet där överträdelsen skett , överträdelsen mot den allmänna ordningen , måste ta sitt ansvar .
Det måste få tillfälle att vidta åtgärder och kommissionen måste upplysas .
Kommissionen måste få möjlighet att kunna agera mot det land som låtit överträdelsen ske .
Grundprincipen i direktivet om elektronisk handel är med andra ord ursprungslandet med en avvikelse som är mycket noga angiven .
Herr talman !
Får jag även ta tillfället i akt att uppmana parlamentet på rätt sätt , det vill säga snabbt , godkänna direktivet så att det kan införlivas i det europeiska rättssystemet efter rådet ( inre marknaden ) i maj i år .
Var och en väntar på ett europeiskt direktiv om elektronisk handel och jag hoppas att vi kan lägga fram ett sådant i maj .
Herr talman !
Jag skulle gärna vilja ta upp ett annat ämne som också nämnts av ett antal parlamentsledamöter .
Inte minst av Palacio men även av Oomen , och det gäller Brysselkonventionen .
Jag inkasserar kritiken från Palacio om det sätt på vilket kommissionens förslag kommit till stånd .
Vi tar lärdom av det .
Jag skulle dock vilja uppmana parlamentet och i synnerhet utskottet för rättsliga frågor och den inre marknaden att bilda sig en uppfattning om den svåra punkten i artikel 15 .
Ser jag rätt , herr talman ?
I så fall avviker nämligen artikel 15 i kommissionens förslag om Brysselkonventionen på en viktig punkt från den ursprungliga konventionen till förmån för konsumentskyddet .
I den ursprungliga konventionen från 1968 ställs ju två villkor för konsumentens möjlighet att åberopa sina egna rättigheter .
Av de två villkoren har ett försvunnit i kommissionens förslag .
Det är en sak som är av stor betydelse och som också lett till oro bland de olika organisationer som engagerar sig i den här saken .
Det är ett ämne som håller kommissionen sysselsatt .
Jag skall själv hålla ett litet sammanträde nästa vecka tillsammans med fyra andra kommissionsledamöter , bland andra kommissionär Byrne , kommissionär Vitorino och kommissionär Liikanen , för att närmare fundera över artikel 15 .
Jag skulle dock samtidigt , om ni tillåter , herr talman , och om Palacio tillåter , utskottet för rättsliga frågor att å sin sida också uppmärksamma artikel 15 så att kommissionen i ett tidigt skede vet vad Palacios utskott anser .
Wallis talade med rätta om begreppet " joined up administration " .
Låt oss nu i samråd med parlamentet komma fram till en noggrannare begreppsdefinition angående artikel 15 enligt definitionen i kommissionens förslag .
Dessutom har ett antal parlamentsledamöter , Wallis , Oomen och naturligtvis även Palacio , talat om å ena sidan small claim procedures och å den andra sidan om alternative dispute settlements .
Parlamentet måste förstå att det inte är några frågor som ligger direkt inom mitt behörighetsområde .
Det är snarare saker för min kollega Vitorino .
Det hindrar inte att det naturligtvis finns ett nära samband med hela den här frågan .
De två påskyndade och förenklade metoderna för att avgöra juridiska tvister hänger naturligtvis också nära samman med den inre marknadens funktion .
Därför känner jag mig själv i hög grad förbunden med det här ärendet .
I ärlighetens namn måste jag dock säga att Antonio Vitorino ändå i första hand är ansvarig för det .
Jag sade nyss att vi , fyra eller fem kommissionärer , skall träffas nästa vecka onsdag .
Jag lovar att jag skall betona och be om uppmärksamhet för nödvändigheten av att komma fram till de två påskyndade och förenklade metoderna för att avgöra små juridiska tvistemål angående e-commerce .
Jag skulle gärna vilja sluta med att upprepa denna lilla anmärkning .
Vi försöker leta efter jämvikten .
Vi försöker hitta en jämvikt .
Vi vill å ena sidan inte ha det som MacCormick sade .
Vi vill inte ha några long distance rip-offs .
Det vill vi inte .
Jag tackar MacCormick för det färgstarka uttrycket .
Å andra sidan vill vi inte heller det som Wallis sade om att ett överdrivet skydd leder till överträdelser av den inre marknaden .
Det vill vi inte .
Vi vill inte det ena men vi vill inte heller det andra .
Vi måste försöka hitta den rätta vägen mellan de olika faror som lurar , till förmån för den inre marknaden , det vill säga : alla konsumenter i Europa .
Jag förklarar debatten avslutad .
 
Kvinnor och vetenskap Nästa punkt på dagordningen är betänkande ( A5-0082 / 1999 ) av McNally för utskottet för kvinnors rättigheter och jämställdhetsfrågor om meddelandet från kommissionen om " Kvinnor och vetenskap " - Berika den europeiska forskningen genom ökat deltagande från kvinnor ( KOM ( 1999 ) 76 - C5-0103 / 1999 - 1999 / 2106 ( COS ) ) .
( DE ) Herr talman !
Jag vill inledningsvis rikta mitt tack till McNally som på grund av brådskande förpliktelser inte kunde närvara för att själv presentera sitt betänkande här i dag .
Kvinnor och vetenskap - mobilisering av kvinnor i den europeiska forskningens intresse .
Meddelandet inriktas mot två mål : Det ena är att stimulera till diskussion medlemsländerna emellan och att understödja de bästa metoderna för att hjälpa fram kvinnor på områdena vetenskap och teknik .
Det andra är att öka antalet kvinnor som deltar i de forskningsuppgifter som backas upp av unionen , varvid hänsyn tas till åtagandena i unionsfördraget om att skapa lika möjligheter för alla och att höja kvalitén på forskningen , dvs. att driva igenom gender mainstreaming .
Området forskning och teknik är trots allt efter jordbruk och strukturfonder det tredje starkaste området i EU-budgeten .
Vi välkomnar kommissionens meddelande och dess mål samt uppmanar medlemsländerna att tillsammans med kommissionen fortsätta att eftersträva jämställdhet och samarbete .
Vi uppmanar kommissionen att plocka fram liknande och bättre fakta på området kvinnor och vetenskap , att dra upp riktlinjer och föreslå ytterligare åtgärder för att om två år lägga fram en särskild rapport för oss här i parlamentet .
Kommissionen fortsätter sitt arbete för bättre jämförelse mellan sakuppgifterna och vetenskapskvinnorna , kommissionen vill anordna möten med relevanta parter liksom sammanföra de nationella tjänstemännen och vetenskapskvinnorna och alla inblandade i två större konferenser .
Föredraganden välkomnar uttryckligen de åtgärder ur femte ramprogrammet för forskning som nu har vidtagits för att öka antalet kvinnor som deltar och kravet på att andelen kvinnor skall ligga på 40 procent såväl när det gäller Marie Curie-stipendierna som i alla rådgivande organ , liksom de åtgärder som redan föreslagits för det sjätte ramprogrammet för forskning .
Den kvinnliga underrepresentationen inom vetenskaplig forskning har en lång tradition , och det har krävts en hård kamp av kvinnorörelsen för att nå dit man har nått .
I början av århundradet fick de första europeiska kvinnorna besöka ett universitet i Finland .
Ändå är universiteten ännu i dag högborgar av manlig dominans .
I dag är nästan hälften av de studerande kvinnor .
I mitt hemland Tyskland var kvinnorna 1995 för första gången i majoritet på grundkurserna .
För alla studerande är det europeiska genomsnittet 103 kvinnor på 100 män .
Tyskland ligger här på jumboplats i EU med 77 kvinnor på 100 män .
Förvisso slutför fler kvinnor än män sina utbildningar , närmare bestämt i förhållandet 110 : 100 .
I Tyskland och på Irland underskrids dessa siffror .
Vid studievalet finner man nu två tredjedelar av de kvinnliga studenterna inom språkvetenskap och humaniora ; för naturvetenskap måste det ges många fler impulser .
Sinnet för det naturvetenskapliga och tekniska måste väckas i föräldrahemmet och stöttas allmänt av utbildningen , i skolan , på dagis , överallt , och här måste man även slå in på nya vägar .
Samundervisning är inte alltid den enda vägen , även en undervisning uppdelad mellan flickor och pojkar kan ge en impuls just i de naturvetenskapliga och tekniska ämnena .
Kvinnors växande kvalifikationer har dock inte slagit igenom på det vetenskapliga området : vid tillsättandet av poster vid högskolorna kan man nu liksom tidigare konstatera att situationen är katastrofal , antalet ordinarie professurer ligger i unionen på 5 procent , det är en obetydlig ökning jämfört med början av 1900-talet .
Kvinnors jämställdhet inom vetenskapen måste dock leda till att kvinnors innehållsliga inflytande ökar .
Kvinnor och genusforskning är att betrakta som grundforskning , vilken är enormt viktig för Europeiska unionen .
Med hjälp av nya instrument som medlemsländerna är tvungna att utveckla måste den outnyttjade potentialen hos alla kvinnor ökas i forskning och undervisning , och utbytet av erfarenheter främjas .
Nätverk av vetenskapskvinnor måste understödjas och innovativa projekt främjas och byggas ut .
Så kan man exempelvis påvisa ett ökat antal kvinnor inom naturvetenskaperna i Spanien och Italien .
Detta måste undersökas mer noggrant .
Exempel kan man finna också i Tyskland : Under Expo 2000 i sommar kommer ett internationellt kvinnouniversitet för teknik och kultur att äga rum under 100 dagar i Hannover .
Tusen blivande vetenskapskvinnor och 100 kvinnliga professorer arbetar där med ett tvärvetenskapligt forskningsorienterat program på sju projektområden : intelligens , information , kropp , vatten , stad , arbete och migration .
Dessa värdefulla erfarenheter måste samordnas och utvärderas noggrant , och sedan måste beslut fattas om huruvida universitetet kan fortsätta drivas som virtuellt campus med hjälp av modern informationsteknik .
Som medgrundare till kvinnouniversitetet är jag övertygad om att denna think tank kan ge en hint om lösningen på många av våra problem .
EU får med tanke på den europeiska forskningen och dess ställning i globaliseringens tecken inte försitta några chanser .
En chans kommer FN-konferensen Peking + 5 att ge vid halvårsskiftet i New York .
Här kommer man att granska resultaten av uppnådda eller också missade mål .
Genom att de politiskt ansvariga i Europeiska unionen , i alla medlemsländer , agerar konsekvent skall vi komma dithän att vi tillsammans med ledningen för högskolorna , med utskotten vid forskningsinstitutionerna liksom med näringslivet kan utföra riktade strukturella förändringar av ramvillkoren och inleda en förvandlingsprocess som skall utföra gemenskapsuppgiften jämställdhet , så som det föreskrivs oss i Amsterdamfördraget .
Vår framtid kommer - som föredraganden McNally så riktigt säger i sin analys - att finnas på 2000-talet .
Det går inte med något slags smink .
Här måste vi skapa djärva vändpunkter .
Än en gång hjärtligt tack till föredraganden McNally !
Herr talman !
Jag vill börja med att klargöra att jag talar för Elisabeth Monforts räkning , vilken är talesman för UEN-gruppen i denna fråga och således kommer jag att läsa den text hon har förberett på franska .
Herr talman , lyckligtvis har det funnits ett brett samförstånd om den debatt som inletts inför utskottet för industrifrågor , utrikeshandel , forskning och energi om betänkandet McNally , i synnerhet i syfte att öka och underlätta kvinnors deltagande i forskningsyrkena .
För att undvika en viss förvirring behöver vi emellertid fördjupa begreppet lika möjligheter som inte verkar omfatta samma verklighet för alla .
I den första versionen av yttrandet hade man bestämt sig för en definition som inte bara var förenlig med kvinnornas legitima ambitioner att få lika tillträde till vetenskapliga studier och att snabbt få medföljande åtgärder som gör det möjligt för dem att få anställningar med ansvar som överensstämmer med deras resultat , men också med begreppet komplementaritet , det enda som kan berättiga en voluntaristisk politik i frågan .
Parlamentets överväganden bör grundas på dessa värden , som respekterar skillnader , och inte på ett postulat om lika möjligheter för kvinnor och män som inom sig bär sina egna motsägelser .
Om nu män och kvinnor är exakt lika och om kvinnan när allt kommer omkring bara är en människa som en annan , finns det inte något skäl för att vilja föreskriva någon jämställdhet mellan kvinnor och män och bara kompetenskriterier bör vara gällande vid fördelningen av tjänster .
Det är således accepterandet av skillnaden och förutfattade meningar om komplementaritet som tvärtom bör återställa balansen och tjäna som stöd för en voluntaristisk , realistisk och pragmatisk politik enligt vilken man framför allt ser till att avskaffa konkreta hinder och de specifika hinder huvudsakligen på grund av förhållandet att de är mödrar , som bara kvinnor har .
En godtycklig kvantitativ politik som vilar på användning av kvoter kommer inte att bidra till att lösa de grundläggande problemen .
Det skulle vara bra om parlamentet gav uttryck åt sin goda vilja rörande kvinnors tillträde till vissa yrken , i synnerhet forskningsyrkena , där de ännu i hög grad är underrepresenterade , i formuleringar som slutgiltigt lägger de retoriskt uttryckta kraven på hyllan .
Herr talman !
Män och kvinnors lika rättigheter regleras i artikel 2 och 3 i Amsterdamfördraget och är därmed ett av de mål som Europeiska unionen alltid skall beakta i sin gemenskapspolitik .
Antalet kvinnor inom det vetenskapliga området har de senaste åren ökat kraftigt , men det räcker inte .
Antalet kvinnor på universitet ökar , på alla områden , men på de utbildningar som vi skulle kunna kalla " vetenskapliga " - som till exempel matematik , data , ingenjörsvetenskap och arkitektur - är de fortfarande underrepresenterade .
Efter avklarade studier med goda betyg fortsätter de inte heller den vetenskapliga utbildningen , mycket på grund av alla hinder som uppstår , vilket förvärrar situationen än mer .
En orsak är upplägget av den vetenskapliga utbildningen och en annan hur de skall kompromissa mellan yrkeslivet och familjelivet .
Därför tycker vi att kommissionens vilja och det intresse man där visar för att försvara kvinnors delaktighet inom vetenskapen , i specifika program , är av stor vikt , även om det mest intressanta för oss är deras delaktighet i det femte ramprogrammet för forskning teknisk utveckling och demonstration ( 1998-2002 ) .
De åtgärder som skall vidtas för att integrera kvinnorna bör finnas med i de särskilda program som tidigare nämnts .
Kvinnan kan med sina speciella egenskaper starkt bidra till forskningen ock kommer utan tvekan att berika vetenskapen .
Ett jämlikt deltagande bör främjas , där målet bör vara jämlikhet , utan att för den skull förglömma att yrkeskunskaper är ett absolut måste .
Kvinnor inom det här området måste gynnas redan på universitetsnivå , särskilt på de mera vetenskapliga utbildningslinjerna , och därefter under hela yrkeskarriären .
Unga kvinnliga forskare bör gynnas medelst Marie Curie-stipendium , så att de får tillräckliga medel .
Kvinnor skall delta vid all rådgivning och vid allt beslutsfattande , inte bara i den vetenskapliga forskningen , målet är ju att berika och komplettera .
Redan från skolåldern skall kvinnor uppmuntras att delta i vetenskapliga aktiviteter , särskilt när det gäller informationsteknik , eftersom det är mycket viktigt även för andra vetenskaper , inte bara inom Europeiska unionen utan också i våra associerade länder och i de områden i underutvecklade länder där unionen genomför olika program .
Kvinnor skall uppmuntras att delta i vetenskapliga program och i den nya tekniken redan från skolåldern .
Större delaktighet inom vetenskapen skall återspegla den betydelse kvinnor spelar på alla sociala områden .
Större delaktighet i femte och sjätte ramprogrammet är ett exempel på jämlikhet mellan män och kvinnor , detta skall åstadkommas genom att göra det lättare för kvinnor att ta sig in i de sektorer som de traditionellt sett har varit underrepresenterade i .
En kompromiss mellan familjeliv med yrkesliv måste nås så att fler kvinnor kan ta sig an ansvarsfulla befattningar .
I parlamentet - särskilt i utskottet för kvinnors rättigheter och jämställdhetsfrågor - kommer vi att fortsätta att arbeta för att nå de grundläggande målen för ett mera likvärdigt samhälle .
Herr talman !
Jag skulle först vilja ge mina komplimanger till Europeiska kommissionen för det initiativ som den har tagit för att mobilisera kvinnorna med målet att få ett större kvinnligt deltagande i vetenskapen och att berika den europeiska forskningen .
Det är ett faktum att det kvinnliga könets representation på området för vetenskaplig forskning och teknik är mycket låg och inte alls motsvarar de framsteg som har gjorts , delvis tack vare den europeiska politiken , på andra områden .
Särskilt då inom utbildningen , där vi verkligen kan tala om en kvinnornas triumf , eftersom kvinnorna på nästan alla europeiska universitet utgör en majoritet av studenterna .
Gröner presenterade tidigare många och intressanta siffror .
Kvinnornas ställning i allmänhet inom den vetenskapliga forskningen med avseende på karriärsplatser hänger naturligtvis i hög grad samman med deras val i utbildningssystemet , men även med deras ställning i familjen .
De olika studieinriktningar som de två könen följer påverkar deras framtida utveckling .
Det är därför nödvändigt att vi i god tid ingriper redan vid yrkesorienteringen i skolan , och att vi informerar de unga kvinnorna om de följder som deras val får för deras yrkesliv .
Å andra sidan påverkar de kvarlevande traditionella rollerna och uppdelningen av arbetet efter kön kvinnornas utveckling och karriär negativt .
Därför är åtgärderna som avser att göra det möjligt att förena familjeliv och yrkeskarriär naturligtvis fortfarande nödvändiga .
Men jag skulle säga att det måste gälla framför allt för männen .
Det är nödvändigt att männen förenar karriären med deltagande i familjelivet , i det privata livet .
Kvinnorna utgör hälften av den mänskliga potentialen , hälften av den globala källan för talang , begåvning och kreativitet .
Att bevara den nuvarande obalansen på det viktiga forskningsområdet är samma sak som att slösa bort värdefulla resurser .
Frågan hör faktiskt samman med Europeiska unionens utveckling och framtid .
Inte en enda av dagens utmaningar kan bemötas utan det bidrag som kvinnornas idéer , fantasi och begåvning utgör .
Utöver kravet på rättvisa mellan de två könen , har alltså frågan också en tillväxtdimension .
Det vill säga nödvändigheten av att stärka konkurrens- och innovationskraften i unionen .
Vad gäller det femte ramprogrammet , har det även som mål att integrera politiken för jämlikhet mellan könen .
Vi stöder de initiativ som mobiliserar kvinnornas många vetenskapliga nätverk och som säkerställer ett könsbalanserat deltagande i de kommittéer och organ som utformar strategier , väljer ut och bedömer projekt och beslutar om vart medlen skall gå .
Vi uppmanar Europeiska kommissionen och medlemsstaterna att undersöka i vilken utsträckning kvinnorna är tillräckligt representerade i den gemensamma jordbrukspolitiken , i strukturfonderna , i det femte ramprogrammet , i de många vetenskapliga och tekniska kommittéerna liksom även i nyckelpositioner .
För att avsluta , herr talman , skulle jag vilja be Europeiska kommissionen att sätta som mål att , genom programmen för föranslutningsstöd till ansökarländerna och till Turkiet , utveckla kvinnornas vetenskapliga talang och att öka kvinnornas möjligheter att bidra till den vetenskapliga och tekniska forskningen och utvecklingen .
Herr talman , kommissionär Busquin , kolleger !
Vi i Gruppen De gröna / Europeiska fria alliansen har läst McNallys betänkande om kvinnor och vetenskap med stort intresse och vi är naturligtvis inte nöjda med den obalans som finns mellan kvinnornas ställning i vetenskapen och männens ställning .
Vi tycker dock att det är viktigt att den här situationen blir belyst och att det läggs fram förslag om en förbättring av kvinnornas ställning .
Kommissionär Busquin har också offentliggjort en rapport angående en studie som gjorts på uppdrag av Europeiska kommissionen .
Tolv kvinnliga vetenskapsmän från olika medlemsstater har tagit fram hårda siffror som visar obalansen i den vetenskapliga världen .
Dessutom har de lagt fram mycket konkreta förslag om förbättring av den nuvarande situationen för kvinnorna .
Av studien framgår också tydligt att orsaken till den här obalansen måste åtgärdas i vetenskapsvärlden i sig och att åtgärderna inte skall beröra kvinnor som skulle ha andra intressen och ambitioner och som skulle göra andra yrkesval .
Det visar sig vara fördomar .
Både i universiteten och i forskningsinstituten och inom industrin så finns det problempunkter .
Inom var och en av dessa arbetskretsar är det på nytt en obalans i fördelningen av funktionerna .
Andelen kvinnliga professorer varierar till exempel i medlemsstaterna från 4 procent till högst 18 procent av hela kåren .
Dessutom visar det sig att andelen kvinnliga professorer i en och samma institution är betydligt mindre än andelen kvinnliga assistenter .
Av en analys av ansökningsuppgifter framgår det att kvinnor som tydligt satsar på en vetenskaplig karriär väljs ut i mycket mindre antal än deras manliga kolleger .
Inte ens barn verkar i det här fallet vara ett hinder , tvärtom , kvinnor med barn och familj skulle till och med publicera mer än ensamstående .
Anmärkningsvärt är att andelen kvinnor med ett vetenskapligt arbete är högre i de sydeuropeiska länderna än i de nordeuropeiska .
En förklaring till det är att det i de senare länderna är lättare att få längre ledigheter men det har också till följd att det inte längre är så självklart att komma tillbaka i den vetenskapliga karriären .
Man bör alltså vara ytterst vaksam när det gäller kvinnor och familjevänliga regler och vidta nödvändiga åtgärder för att kvinnorna verkligen skall få behålla lika möjligheter som männen .
Vi hoppas att den här studien , tillsammans med McNallys betänkande skall vara en ansats till ytterligare initiativ för att fylla upp behovet av siffermaterial .
Vi räknar med att Europeiska kommissionen vidtar åtgärder för att skapa sådana förhållanden att de förslag som lagts fram kan omsättas i praktiken .
Jag skulle vilja avsluta med kommissionär Diamantopoulous ord : vi kämpar för våra rättigheter och inte för några privilegier .
Herr talman , kära kolleger , låt mig bara i första hand säga att jag tycker det är litet synd att debatten om " Peking + 5 " redan sköts upp till slutet av parlamentssammanträdet för en månad sedan , liksom nu på nytt " Kvinnor och vetenskap " .
Så snart det handlar om kvinnor verkar det som att man alltid skjuter upp diskussionen till slutet av alla debatter .
Jag beklagar det .
Herr talman , kära kolleger , när vi läser betänkandet McNally vet vi omedelbart att vi där närmar oss en väsentlig fråga .
" Kvinnor och vetenskap " är en titel som skulle kunna vara bedräglig om man förde in den i en förteckning som för alltid är ofullständig om " Kvinnor och ... " det och det ämnet : en uppräkning är nödvändig men ibland ineffektiv för att förklara ett problems betydelse .
Vi berör här en väsentlig fråga som sedan århundraden tillbaka väcker stridigheter om jämlikheten mellan kvinnor och män .
Kan kvinnor ha samma skäl som män ?
Är kvinnor i stånd att ha en vetenskaplig verksamhet ?
En del tvivlar ännu på det och likväl är svaret hädanefter och för alltid : ja .
Men där börjar svårigheterna .
Om kvinnornas situation på det vetenskapliga området är oroande beror det på en rad problem som är svåra att lösa .
Vetenskap , en symbolisk verksamhet , är ett manligt privilegium , på samma sätt som det politiska ansvaret .
Man finner samma låsningar när det handlar om att dela den politiska makten som när det handlar om makten över tanken .
I båda fallen står den manliga makten på spel .
Låt oss då föreslå samma botemedel , såsom införandet av jämställdhet inom politiken som prövas av vissa länder i unionen .
Flickor lyckas utmärkt i skolan och det finns ingenting som berättigar till att de är så få i forskningsvärlden .
Hindren för en vetenskaplig karriär finns utanför själva forskningen .
Med andra ord räcker det inte att få tillträde till det vetenskapliga området , det måste också finnas plats för kvinnor på området , det vill säga andra kvinnor än de evigt inbjudna , såsom det sades så bra på det möte som hade ordnats av kommissionen i april 1998 .
Studievägledningen inom skola och universitet är en gåta när det gäller jämlikhet mellan kvinnor och män .
De exakta vetenskaperna ordnas ofta på så sätt att de avskräcker flickorna .
Samundervisning liksom eventuell könsdiskriminering av lärare , föräldrar och institutioner är långt ifrån lösta problem .
Vad beträffar de mänskliga vetenskaperna kommer de bara att få en mening om de införlivar kravet att tänka på dimensionen " man-kvinna " i samtliga sociala och mänskliga problem .
Man måste självklart ha en bred vision om vetenskap , och man måste veta att man inte kan tänka ut ett samhälle utan att införa dimensionen " man-kvinna " .
Vi har för närvarande långt kvar .
Jag uppskattar betänkandet McNally för att det är lika fullständigt som sammansatt .
Det verkar viktigt för mig eftersom hon betonar botemedlen , eller rent av lösningarna , i betänkandet för det problem som det svåra utövandet av vetenskap utgör .
Det vill säga hon lämnar i synnerhet uppgifter , naturligtvis med beräkningar , om kvinnornas närvaro inom de olika yrkessektorerna , stipendier och diplom , införandet av tvingande åtgärder för att öka kvinnors närvaro inom forskningen samt främjande av undersökningar om könsdiskrimineringens mekanismer , inrättande av arbetsgrupper och vaktinstanser i kommissionens generaldirektorat Jag gläder mig åt att hon i betänkandet inte har utelämnat vare sig problemet om kvinnors makt inom vetenskapen , ...
( Talmannen avbröt talaren . )
Herr talman !
Kravet på lika villkor för kvinnor och män har visserligen hög prioritet i fördragen , exempelvis i artiklarna 2 och 3 i Amsterdam-fördraget , men i yrkeslivet finns det väsentliga brister .
På området vetenskap och teknik - det aktuella ämnet - finns detta med endast i form av de mest blygsamma ansatser .
Här är kvinnorna snarast sysselsatta i osäkra jobb .
De har lägre inkomster än män .
Inte ens 10 procent är anförtrodda forskningsuppgifter för att inte säga ledarpositioner .
Den låga representationen av kvinnor motsäger absolut deras talanger och förmågor , deras höga nivå av kreativitet och flexibilitet .
Det finns redan i dag europeiska program som lämnar betydande bidrag i syfte att förbättra kvalitén på forskningsresultat , men också att fördjupa samarbetet medlemsstaterna emellan .
En bas för förändringar till det bättre är å ena sidan statistiskt material med könsspecifika fakta och å andra sidan kunskapen om olika modeller för att hjälpa fram kvinnor .
Andra program i gemenskapen , såsom delar av Sokrates och Leonardo för bildning och utbildning , skall överlappas med åtgärder på nationell nivå , såsom läroplaner som i ökad utsträckning innehåller ämnena matematik och naturvetenskap .
Då kommer unga kvinnor att erövra tillgången till informationsteknologin .
Många av dem kommer att bli erkända vetenskapskvinnor .
De kommer alltså att göra karriär , för en gångs skull inte på de klassiskt kvinnliga domänerna , dvs. yrken inom utbildning , medicin eller det sociala .
Vad krävs ?
Fler deltidsarbetsplatser , fler inrättningar för barnomsorg på företagen och alldeles särskilt fler kvinnor i rådgivnings- , urvals- och beslutsorganen för projekt och positioner .
Emellertid kan jag inte helt och hållet dela synen på kvoteringstvång .
Att statiskt låsa sig vid att antalet kvinnor skall vara 40 procent i forskningsprogram och institutioner skadar självförtroendet hos de kvinnor som tagit sig fram eller kommer att ta sig fram utan dylika så kallade hjälpinsatser .
Som en flexibel riktlinje eller som orienteringspunkt kan jag dock absolut acceptera detta med hänsyn till den iögonenfallande underrepresentationen av kvinnor i vetenskapen .
Herr talman !
Jag vill först och främst gratulera kommissionen till lämpligheten och kvaliteten i dess meddelande om kvinnor och vetenskap i vilken påvisas den existerande obalansen och behovet att förändra denna situation .
Jag vill också gratulera min kollega Eryl McNally till det utmärkta betänkandet som hon har utarbetat och till de förslag hon har lagt .
Ur min utgångspunkt kunde detta betänkande inte ha kommit vid ett lämpligare tillfälle .
Det är ett erkänt faktum att kvinnornas deltagande i det aktiva livet är väsentligt för Europas framtid .
Sysselsättningsnivån i Europa är lägre än i USA och Japan , och till detta faktum bidrar den fortfarande låga nivån av kvinnlig medverkan i de flesta av unionens länder .
Om kvinnors roll är viktig för att öka den europeiska produktionen , är betydelsen av deras bidrag till finansieringen av social trygghet och alltså bibehållandet av en social modell , också värt att nämna .
Men det räcker inte med att analysera kvantiteten arbete som utförs av kvinnor i Europeiska unionen .
För oss är också det utförda arbetets kvalitet och samhällets erkännande av stor vikt vilka , sammanbundna med kvinnornas professionella kvalifikationer , måste ligga i nivå med deras närvaro i de mest krävande branscherna vad gäller yrkesutbildning och där ligger Europeiska unionen mycket långt efter .
I Europeiska unionen finns i själva verket mellan 700 000 och 800 000 lediga platser på grund av brist på rätt utbildad personal för att utveckla informationssamhället och användandet av nya tekniker .
Vetenskapskvinnorna i Europa måste alltså ges allt stöd och öppningar för att de skall få sin rättmätiga roll vilket Europa också är i behov av .
Jag knyter tidpunkten för detta betänkande till att det portugisiska ordförandeskapet skall genomföra ett extra toppmöte i Lissabon i mars , om sysselsättning , ekonomiska reformer och sammanhållning för ett Europa med innovation och kunskap , vilket skall försöka skapa grunden för en utvecklingsmodell som placerar Europa i täten för den ekonomiska konkurrenskraften på internationell nivå .
Detta är inte möjligt utan ett enormt deltagande från de vetenskapskvinnorna i Europa .
Därför måste vi sätta in positiva åtgärder i denna fråga och inte bara låta utvecklingen av ett samhälle och en politik som är mer mainstream ske av sig själv .
Jag har välgrundade förhoppningar om att det portugisiska ordförandeskapet skall uppmärksamma kvinnornas medverkan i detta program på vederbörligt sätt , inte bara därför att det portugisiska Jämställdhetsministeriet är knutet till det , utan också för att den portugisiske premiärministern - och inte av en slump - gav samordningen av det program som skall läggas fram på toppmötet i Lissabon i uppgift till en vetenskapskvinna .
Jag hoppas att kommissionens och rådets goda intentioner resulterar i konkreta förslag för att få ett större deltagande av de europeiska kvinnorna , kvantitativt och kvalitativt , på de vetenskapliga och de nya teknikområdena .
Herr talman , kolleger !
Vi undersöker i dag problemet med kvinnornas tillträde till vetenskap och forskning .
Kommissionens text , men även betänkandet , når inte sitt mål .
Till att börja med kopplar de inte ihop ämnet med den mer allmänna kvinnofrågan .
De presenterar inte kvantitativa siffror som skulle ge en tydlig bild av situationen , förutom viss statistik om proportionen mellan könen i universitetsstudierna .
Mellan universitetsstudierna och forskningssysslan är det dock en enormt avstånd .
Det största felet med texterna är emellertid att man inte fördjupar sig i frågan och att de inte pekar på orsakerna till problemen .
Den luddiga hänvisningen till förekomsten av komplexa strukturella barriärer eller till och med till att den rådande mentaliteten på forskningsområdet i allmänhet är maskulin , kan väl inte anses vara allvarliga försök att tolka situationen .
Oförmågan att utveckla produktionsfaktorerna , framför allt den mänskliga , liksom bristen på lika möjligheter , är grundläggande kännetecken för det kapitalistiska systemet .
Det har allvarliga följder för särskilt de känsligaste sociala skikten , dit unga och kvinnor räknas .
Det är ingen tillfällighet att kvinnornas situation och sociala ställning var mycket bättre i de före detta socialistiska staterna än i väst .
Det samhälle som vi lever i har skapat en ram som är fientlig mot kvinnorna .
Till exempel får politiken med ständiga och allt större nedskärningar av välfärden och demolering av de offentliga socialförsäkringssystemen till följd att kvinnan utsätts för ett större tryck att ägna sig åt sin traditionella roll .
Det gäller i högsta grad för kvinnliga forskare .
Helt klart är att problemet inte kan lösas med den så kallade flexibiliteten , inte heller med deltidssysselsättning , eftersom det inte går att bedriva forskning utan att lägga ned mycket tid och arbete .
Mot många av förslagen i resolutionen , som förslagen om en mer detaljerad statistik , en databas för kvinnliga experter , med flera , finns det knappast någon som har invändningar .
Men problemet kan inte lösas med dessa åtgärder .
Och ännu mindre kan man lösa problemet med kvoter .
Det krävs en annan politik som innebär att människan i allmänhet och kvinnorna i synnerhet respekteras och som inte har fåtalets vinst som drivande kraft och exploateringen av flertalet som mål .
Naturligtvis förväntar vi oss inte att Europeiska unionen skall driva en sådan politik .
Vi förväntar oss dock av folken i Europeiska unionen tvingar fram den .
Herr talman !
Det gläder mig mycket att kunna ta till orda för att meddela att jag stöder programmet som lagts fram av McNally för att ge kvinnorna bättre möjligheter att berika det vetenskapliga området .
För första gången talar jag nu som företrädare för Pensionärspartiet .
Jag är visserligen nationell sekreterare för Pensionärspartiet i Italien , men ordföranden är en kvinna , Giuseppina Cardazzi , och vi inser med andra ord verkligen kvinnornas betydelse .
Inom inget annat område är det lika viktigt som inom forskningen att man förverkligar jämlikheten mellan män och kvinnor .
Hittills har vi haft - för att bara nämna ett par exempel - enbart manliga vetenskapsmän , som Leonardo da Vinci , Michelangelo , von Braun , Einstein etc .
Föreställ er , kommissionär Busquin , att kvinnorna under de senaste två tusen åren hade haft samma möjligheter som männen !
Föreställer er , herr talman , om kvinnorna sedan två tusen år tillbaka hade befunnit sig i den situation dit kommissionen vill föra dem i och med detta förslag .
Jag är helt övertygad om att om det hade varit på det viset , så hade vi i detta ögonblick kommit betydligt längre i vår utveckling än vad som nu är fallet .
Kvinnorna lever som bekant betydligt längre än männen .
Vi frågar oss vad det är de har utöver det som männen har , men jag är övertygad om att detta något , som vi ännu inte känner till , kommer att visa sig även inom den vetenskapliga forskningen .
Förslaget blir desto viktigare som det tillåter kvinnorna att utveckla denna sin vetenskapliga kapacitet - som hittills har legat dold - snarare än att det erbjuder dem arbetstillfällen .
Därför är jag speciellt lycklig över att kunna ge mitt stöd till detta betänkande .
Herr talman , mina damer och herrar !
Av erfarenhet vet vi att den som inte talar om sig själv tyvärr ofta glöms bort , och det är vad vi diskuterar i kväll .
Tusen tack , herr kollega , för de vänliga , uppmuntrande orden .
Men av erfarenhet , och av talen som har hållits här i kväll , vet vi ju också att det inte är den goda viljan det hänger på och inte heller på kvinnorna själva .
Det är ett komplext , strukturellt motstånd , ja man skulle kanske också kunna säga ett kvinnotypiskt motstånd , som har gjort att det fortfarande inte är möjligt för kvinnor att i högre grad vara aktiva inom vetenskap och forskning .
Här är vi kvinnor underrepresenterade , och ingen av talarna här i kväll har heller påstått något annat .
Vetenskap och forskning - den som vill arbeta inom detta område , den som vill ha möjligheter här , han eller hon måste också kontinuerligt kunna avancera .
Och även det är ofta ganska så , ganska så svårt för kvinnor .
Man måste vara flexibel .
Kvinnor är bundna till familj , barn , kanske även till makens arbetsplats .
Då måste man erbjuda flexibilitet , gå kvinnorna till mötes och sedan också ge dem möjlighet till en kontinuerlig vidareutveckling på detta så rasande snabba område .
Det femte ramprogrammet arbetar i synnerhet på att inbegripa frågan om lika möjligheter .
EU : s förpliktelser i fråga om jämställdhet måste ge utslag alldeles särskilt på det vetenskapliga området .
Instrument och metoder för att ge handledning i de klassiska naturvetenskapliga ämnena redan åt flickor måste helt enkelt också få stöd .
Kvinnor bevisar sin akademiska förmåga på de vetenskapliga utbildningslinjerna , och likafullt får vetenskapskvinnorna ännu i dag lägre lön än sina manliga kolleger .
De innehar sällan en ledande position , står sällan i ansvarsställning .
Vetenskaplig forskning som gjorts av en kvinna respekteras ofta mindre än de manliga kollegernas forskning utav expertkommittéer .
Vi har nått enighet här i detta rum i kväll .
Vi gläds åt kommissionsrapporten och hoppas att vi därmed också skall göra framsteg på vägen mot fler kvinnor inom vetenskapen . )
Principen om lika rättigheter betraktas som fundamental och genomsyrar all gemenskapspolitik , vetenskapen får inte vara ett undantag .
Därför måste vi välkomna McNallybetänkandet samt därtill hörande uttalande från kommissionen med den förhoppningen att kammaren ger den sitt fullständiga stöd .
Jag vill ta upp tre frågor som jag anser vara av särskilt intresse .
Den första åsyftar , precis som det påpekas i betänkandet och i uttalandet , att det är länderna i söder - Italien , Portugal och Spanien - där kvinnans närvaro på det vetenskapliga området är mera jämställd , vilket visar att det är viktigt , som i det dagliga livet , att inte tro på alla klichéer .
Den andra frågan berör kvoterna .
Det är omöjligt att inte beakta kvantitativa faktorer vid utvärderingen av en politik , men kvoterna måste tolkas mera allmänt för att se vilka tendenser som finns , det vill säga som ett mål som vi på kort eller längre sikt bör nå , något vi bör tillämpa i mera allmänna ordalag och inte som en siffra som vi hårdnackat och automatiskt måste ålägga varje rådgivande grupp och varje utvärderingsgrupp .
Incitament , stimulans , befrämjande åtgärder , eliminering av hinder och annat som kan vara till förfång måste utan avbrott försöka åstadkommas .
Vad vi i alla fall aldrig kan göra är att spänna spannet före oxarna .
Det är det gamla problemet om mål och medel .
Medlen måste vara lämpliga och väl avvägda och de får framför allt inte äventyra det högsta goda , det vill säga kvalitet , rigorism och räckvidd inom vetenskapen .
Avslutningsvis så är den tredje frågan den att vetenskapliga metoder inte har något kön .
Madame Curie tänkte på samma sätt som Lord Rutherford och madame Kowaleska tänkte på samma sätt som Elie Cartán .
Vi måste göra allt som står i vår makt för att öka kvinnors närvaro inom vetenskapen , men låt oss inte ta en genväg så att vi tappar bort oss .
( Applåder ) .
( FR ) Herr talman , när kommissionen lade fram meddelandet ville den ta ett starkt politiskt initiativ i frågan om kvinnornas plats inom forskningen .
Jag gläder mig åt att konstatera att initiativet har tagits emot väl av parlamentet , som jag tackar för den viktiga roll som det spelar i dynamiken " kvinnor och vetenskap " .
Det resolutionsförslag som vi diskuterar i dag stöder i stort de riktlinjer som kommissionen utarbetat .
Det är en stor och betydelsefull uppmuntran .
Men frågan om kvinnor och vetenskap ingår i ett bredare perspektiv om unionens forskningspolitik .
Såsom jag redan angav till utskottet för industrifrågor , utrikeshandel , forskning och energi är målet att utveckla en politisk strategi för att skapa ett europeiskt område för forskning .
Kommissionen har just godkänt ett meddelande i det avseendet den 18 januari .
Inrättandet av ett sådant område kommer att göra det möjligt att bättre mobilisera den potential vetenskapskvinnorna utgör och att anta den gemensamma utmaningen rörande kvinnors underrepresentation inom forskningen .
Kommissionen är medveten om debatten om principen om kvoter på området för kvinnors deltagande i allmänhet .
Denna debatt utökas naturligtvis till att röra kvinnors deltagande i vetenskaplig forskning .
Kommissionen har inte valt angreppssättet med obligatoriska kvoter utan föredrar kvantitativa mål för deltagande tillsammans med en uppföljning och en utvärdering .
Kommissionen anser att med detta angreppssätt kan man få kvinnors deltagande att öka samtidigt som man respekterar principen om vetenskaplig högsta kompetens .
Betänkandet McNally , som enhälligt godkändes av utskottet för kvinnors rättigheter och jämställdhetsfrågor , stöder kommissionens riktlinjer , vars mål är att uppnå minst 40 procent kvinnligt deltagande i vissa delar av genomförandet av det femte ramprogrammet .
Detta stöd är viktigt .
Redan nu är kvinnornas närvaro 26 procent i de rådgivande grupperna och 24 procent i kontroll- och utvärderingspanelen , vilket är en avsevärd framgång jämfört med det fjärde ramprogrammet .
Det finns fortfarande ansträngningar att göra , men jag tror att vi har slagit in på rätt väg .
McNally rekommenderar också att undersökningar om genuseffekter i de specifika programmen i det femte ramprogrammet beaktas i det sjätte ramprogrammet .
Anbudsinfordran rörande dessa undersökningar har redan offentliggjorts av kommissionen .
Den sköter utvärderingen av mottagna anbud .
Resultatet av dessa undersökningar kommer att göra det möjligt att fastställa det sjätte ramprogrammets riktlinjer .
Men främjandet av lika möjligheter går längre än den begränsade ramen för gemenskapsprogrammen för forskning och jag förstår att parlamentet är angeläget om att se denna fråga beaktas i unionens övriga politik .
Kommissionen agerar redan inom det området och kommer att fortsätta att göra det .
Till exempel , inom ramen för riktlinjerna för sysselsättningen , den fjärde axeln och i förordningsbestämmelserna rörande strukturfonderna .
I sitt förslag till reform som är föremål för en vitbok sätter kommissionen upp målet om en bred balans när det gäller kvinnors och mäns närvaro på alla områden och på alla tjänstenivåer .
McNally föreslår att vi undersöker orsakerna till att det finns klyftor mellan antalet kvinnor med examina inom de vetenskapliga grenarna och antalet kvinnor som in fine utövade ett yrke på området .
Ett antal talare tog upp denna tanke .
Orsakerna till klyftan är komplexa och den rapport som nyligen publicerades av ETAM : s experter tar upp frågan .
Det är viktigt att vi fortsätter att fördjupa analysen för att bättre identifiera hindren och botemedlen .
I det avseendet fortsätter man för övrigt aktivt med genomförandet av den handlingsplan som lades fram i meddelandet och ETAM : s expertrapport , som Sorensen så relevant har åberopat , gör en sammanfattning av kvinnornas underrepresentation inom forskningen .
Rapporten lades fram den 23 november i närvaro av parlamentsledamöter , bland vilka McNally ingick .
Rapporten som utarbetats av oberoende experter är ett mycket nyttigt instrument för att främja diskussion och klarlägga konkreta åtgärder .
Den slutliga versionen av dokumentet kommer att vidarebefordras till parlamentet .
Men det finns andra utarbetningar på gång .
Jag vill påminna om att i juli ordnades ett sammanträde om vetenskapskvinnors nätverk och en grupp nationella tjänstemän samlades den 29 och 30 november för att jämföra politiska åtgärder för att främja kvinnor på det vetenskapliga området på de olika medlemsstaternas nivå .
I det avseendet vidtar kommissionen åtgärder i samarbete med medlemsstaterna - Gröner har betonat den tyska ansträngningen i frågan i det avseendet .
Med grupper av nationella experter utarbetar vi statistiska indikatorer om kvinnors deltagande i europeisk forskning , eftersom det är mycket viktigt att förfoga över pålitliga indikatorer på alla nivåer och de nationella experterna är i det avseendet mycket nyttiga .
Jag skulle till slut vilja meddela er att det kommer att bli en stor europeisk konferens i Bryssel den 3 och 4 april för att göra en sammanfattning av läget med samtliga berörda parter : nationella parlament , nationella förvaltningar , forskningsinstitut och nätverk .
Ni är naturligtvis mer än någonsin inbjudna att delta i arbetet .
Jag skulle också vilja säga att i enlighet med åtagandena i meddelandet ämnar kommissionen regelbundet informera parlamentet om de uppnådda framstegen .
Såsom ni underströk kommer vi för övrigt att få ett meddelande år 2001 på grundval av samtliga rapporter som utarbetats .
Jag slutar med att säga att frågan " Kvinnor och vetenskap " tvingar oss att se längre än de rena forskningsprogrammen i unionen och bör bli föremål för en bred debatt .
Vi har haft det här , men jag tror och jag skulle vilja tacka er för det , att parlamentets resolution kommer att vara ett betydande stöd i det sammanhanget .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum under nästa sammanträdesperiod .
( Sammanträdet avslutades kl .
20.00 . )
