 
Återupptagande av sessionen Jag förklarar Europaparlamentets session återupptagen efter avbrottet den 17 december .
Jag vill på nytt önska er ett gott nytt år och jag hoppas att ni haft en trevlig semester .
Som ni kunnat konstatera ägde " den stora år 2000-buggen " aldrig rum .
Däremot har invånarna i ett antal av våra medlemsländer drabbats av naturkatastrofer som verkligen varit förskräckliga .
Ni har begärt en debatt i ämnet under sammanträdesperiodens kommande dagar .
Till dess vill jag att vi , som ett antal kolleger begärt , håller en tyst minut för offren för bl.a. stormarna i de länder i Europeiska unionen som drabbats .
Jag ber er resa er för en tyst minut .
( Parlamentet höll en tyst minut . )
Fru talman !
Det gäller en ordningsfråga .
Ni känner till från media att det skett en rad bombexplosioner och mord i Sri Lanka .
En av de personer som mycket nyligen mördades i Sri Lanka var Kumar Ponnambalam , som besökte Europaparlamentet för bara några månader sedan .
Skulle det vara möjligt för er , fru talman , att skriva ett brev till den srilankesiska presidenten i vilket parlamentets beklagande uttrycks över hans och de övriga brutala dödsfallen i Sri Lanka och uppmanar henne att göra allt som står i hennes makt för att få en fredlig lösning på en mycket komplicerad situation ?
Ja , herr Evans , jag tror att ett initiativ i den riktning ni just föreslagit skulle vara mycket lämpligt .
Om kammaren instämmer skall jag göra som herr Evans föreslagit .
Fru talman !
Det gäller en ordningsfråga .
Jag skulle vilja ha råd från er vad gäller artikel 143 om avvisning av ett ärende som otillåtligt .
Min fråga har att göra med något som kommer att behandlas på torsdag och som jag då kommer att ta upp igen .
Cunhas betänkande om de fleråriga utvecklingsprogrammen behandlas i parlamentet på torsdag och det innehåller ett förslag i punkt 6 om att något slag av kvoteringspåföljder bör införas för länder som misslyckas med att uppfylla sina årliga mål rörande minskning av flottorna .
I betänkandet står det att detta bör göras trots principen om relativ stabilitet .
Jag anser att principen om relativ stabilitet är en grundläggande rättsprincip inom den gemensamma fiskeripolitiken , och ett förslag som skulle undergräva den måste betraktas som rättsligt otillåtligt .
Jag vill veta om jag kan göra en sådan invändning mot ett betänkande , som alltså inte är ett lagförslag , och om det är något som jag har behörighet att göra på torsdag .
Det är faktiskt just vid det tillfället som ni , om ni vill , kan ta upp denna fråga , dvs. på torsdag innan betänkandet läggs fram .
Fru talman !
Under årets första sammanträdesperiod för Europaparlamentet bestämde man dessvärre i Texas i USA att nästa torsdag avrätta en dödsdömd , en ung man på 34 år som vi kan kalla Hicks .
På uppmaning av en fransk parlamentsledamot , Zimeray , har redan en framställning gjorts , undertecknad av många , bland annat jag själv , men jag uppmanar er , i enlighet med de riktlinjer som Europaparlamentet och hela den europeiska gemenskapen alltid har hållit fast vid , att med all den tyngd ni har i kraft av ert ämbete och den institution ni företräder , uppmana Texas guvernör , Bush , att uppskjuta verkställigheten och att benåda den dömde .
Detta är helt i linje med de principer som vi alltid har hävdat .
Tack , herr Segni , det skall jag gärna göra .
Det ligger faktiskt helt i linje med de ståndpunkter vårt parlament alltid antagit .
Fru talman !
Jag vill fästa er uppmärksamhet vid ett fall som parlamentet vid upprepade tillfällen har befattat sig med .
Det gäller fallet Alexander Nikitin .
Alla gläder vi oss åt att domstolen har friat honom och tydligt visat att tillgängligheten till miljöinformation är en konstitutionell rättighet även i Ryssland .
Nu är det emellertid så att han skall åtalas på nytt i och med att allmänne åklagaren överklagar .
Vi är medvetna om , vilket vi också - inte minst under förra årets sista plenarsammanträde - har kunnat konstatera i en lång rad beslut , att detta inte enbart är ett juridiskt fall och att det är fel att beskylla Alexander Nikitin för kriminalitet och förräderi , eftersom vi som berörda parter drar nytta av de resultat han har kommit fram till .
Resultaten utgör grunden för de europeiska programmen för skydd av Barents hav , och därför ber jag er granska ett utkast till ett brev som skildrar de viktigaste fakta samt att i enlighet med parlamentsbesluten visa Ryssland denna ståndpunkt klart och tydligt .
Ja , fru Schroedter , jag skall mycket gärna granska fakta rörande denna fråga när jag fått ert brev .
Fru talman !
Först skulle jag vilja ge er en komplimang för det faktum att ni hållit ert ord och att det nu , under det nya årets första sammanträdesperiod , faktiskt har skett en kraftig utökning av antalet TV-kanaler på våra rum .
Men , fru talman , det som jag bad om har inte inträffat .
Det finns nu visserligen två finska kanaler och en portugisisk , men det finns fortfarande ingen nederländsk kanal .
Jag bad er om en nederländsk kanal , eftersom nederländare också gärna vill ta del av nyheterna varje månad då vi blir förvisade till den här platsen .
Jag skulle således på nytt vilja be er att ombesörja att vi också får en nederländsk kanal .
Fru Plooij-van Gorsel !
Jag kan tala om för er att frågan finns på föredragningslistan för kvestorernas möte på onsdag .
Jag hoppas att den kommer att granskas i en positiv anda .
Fru talman !
Kan ni berätta för mig varför detta parlament inte följer den arbetsskyddslagstiftning det faktiskt antar ?
Varför har det inte genomförts något luftkvalitetstest i denna byggnad efter denna mandatperiods början ?
Varför har inte arbetsskyddskommittén haft några sammanträden sedan 1998 ?
Varför har det inte skett några brandövningar i parlamentets byggnader i Bryssel eller Strasbourg ?
Varför finns det inga instruktioner om hur man skall bete sig om det börjar brinna ?
Varför har inte trapporna byggts om efter den olycka jag råkade ut för ?
Varför upprätthåller man inte bestämmelserna om rökfria områden ?
Jag tycker det är skrämmande att vi antar lagstiftning som vi inte själva följer .
( Applåder ) Fru Lynne !
Ni har helt rätt och jag skall kontrollera om allt detta faktiskt inte har gjorts .
Jag skall också överlämna problemet till kvestorerna och jag är övertygad om att de är måna om att se till att vi respekterar de regler som vi faktiskt röstat fram .
Fru talman !
Díez González och jag har ställt några frågor angående vissa av vice ordförande de Palacios åsikter som återgavs i en spansk dagstidning .
De ansvariga har inte tagit med dessa frågor på föredragningslistan , eftersom man ansåg att dessa hade besvarats vid ett tidigare sammanträde .
Jag ber att man omprövar det beslutet , eftersom så inte är fallet .
De frågor som tidigare besvarats handlade om de Palacios inblandning i ett särskilt ärende , inte om de uttalanden som återgavs i dagstidningen ABC den 18 november i fjol .
Kära kollega !
Vi skall kontrollera allt detta .
Jag erkänner att för närvarande förefaller saker och ting litet oklara .
Vi skall alltså se över detta mycket noga så allt blir i sin ordning .
Fru talman !
Jag vill veta om det kommer att gå ut ett tydligt budskap från parlamentet under veckan om vårt missnöje rörande dagens beslut om att vägra en förnyelse av vapenembargot mot Indonesien , med hänsyn till att det stora flertalet i detta parlament har stött vapenembargot mot Indonesien ?
Dagens beslut att inte förnya embargot är oerhört farligt med hänsyn till situationen där .
Parlamentet bör alltså sända ut ett budskap , eftersom detta är vad det stora flertalet vill .
Det är oansvarigt av EU : s medlemsstater att vägra att förnya embargot .
Som olika personer har sagt , är situationen där oerhört turbulent .
Det finns faktiskt en risk för en framtida militärkupp .
Vi vet inte vad som händer .
Så varför skall vapentillverkarna i EU profitera på oskyldiga människors bekostnad ?
( Applåder ) I vilket fall som helst är frågan för närvarande inte föremål för någon begäran om brådskande förfarande på torsdag .
 
Arbetsplan Nästa punkt på föredragningslistan är fastställande av arbetsplanen .
Det slutgiltiga förslaget till föredragningslista som utarbetats av talmanskonferensen vid sammanträdet den 13 januari i enlighet med artikel 110 i arbetsordningen har delats ut .
För måndag och tisdag har inga ändringar föreslagits .
Beträffande onsdag : Den socialistiska gruppen har begärt att ett uttalande från kommissionen om dess strategiska mål för de fem kommande åren samt om kommissionens administrativa reform skall tas upp .
Jag skulle vilja att Barón Crespo , som lämnat begäran , uttalar sig för att motivera den , om han vill , naturligtvis .
Sedan gör vi som vi brukar : vi lyssnar till en talare för och en talare emot .
Fru talman !
Framläggandet av kommission Prodis politiska program för hela mandatperioden bottnar i ett förslag från Europeiska socialdemokratiska partiets grupp som antogs med enhällighet på talmanskonferensen i september samt ett tydligt godkännande från ordförande Prodi som upprepade detta åtagande i sitt anförande i samband med tillträdandet av sitt ämbete .
Detta åtagande är viktigt , med tanke på att kommissionen är det organ som enligt fördragen har ensam initiativrätt , och det utgör därför grunden till parlamentets politiska och lagstiftande verksamhet de kommande fem åren .
Jag vill dessutom , fru talman , påminna om att parlamentet vid två tillfällen under föregående mandatperiod röstade om förtroendet för ordförande Prodi ; man röstade på nytt om detta under denna mandatperiod i juli , och sedan , när den nya kommissionen hade påbörjat sitt arbete , gav man i september en förtroenderöst till hela kommissionen .
Därför har det funnits tillräckligt mycket tid för kommissionen att förbereda sitt program och för att oss att ta del av detta och redogöra för detta inför medborgarna .
Jag vill också påminna om resolutionen av den 15 september , där man rekommenderade att förslaget skulle läggas fram så snart som möjligt .
Det som hände förra veckan - något som inleddes utanför talmanskonferensen , en konferens som endast utnyttjades för att bestyrka och bekräfta det beslut som fattats utanför ramarna för denna - utgör ett dilemma : antingen är det så att kommissionen inte är i stånd att presentera programmet ( i sådant fall bör den klargöra detta .
Enligt ordförandens uttalanden kan man presentera programmet .
Med tanke på att kommissionen företräds av vice ordförande de Palacio , anser jag att vi innan omröstningen sker bör få veta huruvida kommissionen är beredd att lägga fram programmet , så som man kommit överens om ) ; annars är parlamentet inte i stånd att granska programmet , så som vissa tycks anse .
Enligt min uppfattning skulle den sistnämnda hypotesen innebära att vi försummade vårt ansvar som parlament , förutom att man då skulle införa en grundtes , en okänd metod som innebär att de politiska grupperna skriftligen får ta del av kommissionens tankar kring programmet en vecka i förväg i stället för en dag i förväg , som man kommit överens om .
Då bör man tänka på att lagstiftningsprogrammet skall debatteras i februari , och därför skulle vi lika gärna kunna avstå från den debatten , för pressen och Internet skulle redan dagen därpå tillkännage programmet för alla medborgare , och det skulle inte längre finnas någon anledning för parlamentet att ägna sig åt frågan .
Eftersom min grupp anser att parlamentet är till för att lyssna , för att debattera och för att reflektera , anser vi att det inte finns något som rättfärdigar en senareläggning av debatten , och om kommissionen är beredd till det , menar vi att det fortfarande är möjligt att återupprätta det ursprungliga avtalet mellan parlamentet och kommissionen och agera på ett ansvarsfullt sätt gentemot våra medborgare .
Därför innebär förslaget från Europeiska socialdemokratiska partiets grupp , som fru talmannen nämnde , att kommission Prodis lagstiftningsprogram läggs fram på onsdag som planerat , och att man inbegriper förslaget om en administrativ reform , för i annat fall kan en paradoxal situation uppstå : å ena sidan vägras kommissionens ordförande , med ursäkten att det inte finns något dokument , rätten att tala i parlamentet , å andra sidan omöjliggörs en debatt om reformen , eftersom parlamentet inte tidigare har fått ta del av dokumenten i fråga .
Därför ber jag , fru talman , att ni uppmanar kommissionen att uttala sig och att vi därefter går till omröstning .
( Applåder från PSE ) Fru talman , ärade kolleger !
Jag måste säga att jag är något förvånad över kollegan Barón Crespos agerande när han nu kräver att denna punkt på föredragningslistan flyttas till onsdagen .
Herr Barón Crespo !
Ni kunde inte närvara vid talmanskonferensen förra torsdagen .
Det tänker jag inte kritisera : det händer alltid att man har en ställföreträdare .
Kollegan Hänsch var där och företrädde er .
Vi förde en grundlig debatt på talmanskonferensen .
Det var bara er egen grupp som förespråkade det ni nu talar om .
Därefter röstade vi .
Varje ordförande har ju lika många röster som hans eller hennes grupp har medlemmar .
Det röstades på denna punkt .
Omröstningen resulterade vad jag kan minnas i följande siffror : 422 röster mot 180 , med några få nedlagda röster .
Detta betyder att alla grupper , med undantag för de grupplösa - men de är ju heller ingen grupp - var överens , och endast er grupp ansåg att man borde förfara på det sätt som ni har föreslagit här .
Alla andra var av en annan åsikt .
Sådant blev beslutet .
Nu vill jag själv säga något i ämnet .
Vi hyser förtroende för kommissionen , för Romano Prodi , och en mycket stor majoritet av vår grupp uttalade sitt förtroende för Romano Prodi och kommissionen efter en , som alla vet , svår process .
Men vi anser också att vi måste föra en debatt om kommissionens strategi under ordnade former , inte bara utifrån ett muntligt uttalande här i Europaparlamentet utan också från ett dokument som kommissionen har beslutat om och som beskriver programmet för fem år framöver .
Något sådant dokument existerar inte !
( Applåder ) I februari skall kommissionen lägga fram programmet för år 2000 .
Vi har sagt att detta går för sig , om kommissionen inte vill göra klart program 2000 redan i januari , då gör vi det i februari .
Det har vi sagt ja till .
Vi vill ju för den delen inte gräla med kommissionen utan anser att kommission och parlament så långt det är möjligt skall gå samma väg .
Men samtidigt är vi som parlament kontrollinstans gentemot kommissionen .
Och allt som kommer från kommissionen behöver inte nödvändigtvis vara vår åsikt .
Jag vill att vi inom grupperna skall kunna förbereda oss på ett klokt sätt inför en debatt om femårsprogrammet .
Man kan inte förbereda sig genom att sitta här och lyssna på ett uttalande utan att alls veta vad som ligger bakom ett sådant uttalande .
Därför rekommenderar vi - och jag har intrycket att kommissionen likaledes är öppen för den tanken - att debatten om kommissionens långsiktiga arbete fram till år 2000 förs nu i februari - jag hoppas också att kommissionen till dess har kommit överens om ett program att föreslå - och att vi samtidigt i februari kan debattera kommissionens lagstiftningsprogram för år 2000 .
Det är sålunda även av förnuftiga och sakliga skäl som vi bör debattera bägge programmen samtidigt .
Därför tillbakavisar min grupp å det bestämdaste den socialistiska gruppens förslag !
( Applåder från PPE-DE-gruppen ) Fru talman !
Jag vill i första hand klargöra att kommissionen hyser den största respekt för parlamentets beslut , och därmed även för beslutet om fastställandet av arbetsplanen .
Vi respekterar således i det avseendet parlamentets beslut .
Samtidigt vill jag klargöra att ordförande Prodi har lovat parlamentet ytterligare en debatt , precis som Barón påpekade , förutom den årliga debatten om kommissionens lagstiftningsprogram , en debatt om de viktigaste handlingslinjerna under den kommande femårsperioden , det vill säga under denna mandatperiod .
Det jag vill säga , fru talman , är att man i den överenskommelse som uppnåddes i september , gjorde en åtskillnad mellan den debatten och framställandet av kommissionens årliga lagstiftningsprogram .
Och jag vill också , fru talman , säga att vi från kommissionens sida är förberedda och färdiga för denna debatt när än det må vara , att vi är redo att hålla debatten denna vecka , så som man i princip avtalade , med tanke på att utkastet redan har presenterats i ett anförande inför de parlamentariska grupperna .
Därför , fru talman , vill jag än en gång påpeka att vi för vår del har diskuterat igenom åtgärdsprogrammet för de kommande fem åren , och att vi är redo att , när som helst då parlamentet beslutar det , - den här veckan om man bestämmer sig för det - komma och presentera programmet för de kommande fem åren , och sedan nästa månad , programmet för år 2000 , precis som avtalat .
Jag föreslår att vi röstar om begäran från den socialistiska gruppen att på nytt föra upp kommissionens uttalande om dess strategiska mål på föredragningslistan .
( Parlamentet avslog begäran . )
Talmannen .
Beträffande onsdagen har jag också mottagit ett annat förslag beträffande den muntliga frågan om kapitalskatt .
PPE-DE-gruppen begär att denna punkt skall strykas från föredragningslistan .
Vill någon kollega begära ordet för gruppens räkning och motivera denna begäran ?
Fru talman !
Eftersom jag hör att det skrattas bland socialisterna : man har sagt mig att även vida kretsar inom den socialistiska gruppen gärna vill se den här punkten avförd från föredragningslistan , eftersom det vid omröstningen på talmanskonferensen saknades votum för berörda kolleger i den socialistiska arbetsgruppen .
Jag vet inte huruvida denna information stämmer , men vi i PPE-DE-gruppen vore i alla fall tacksamma ifall punkten ströks , då ju parlamentet redan har befattat sig med frågan flera gånger .
Det finns också beslut fattade mot en sådan skatt .
Därför yrkar min grupp på att punkten avförs från föredragningslistan .
Tack , herr Poettering .
Vi skall nu lyssna till Wurtz som skall uttala sig emot denna begäran .
Fru talman !
Jag skulle till att börja med vilja understryka Poetterings bristande logik .
Han har just läxat upp den socialistiska gruppen för att den ändrat sig när det gäller ett beslut som fattats med mycket liten marginal i talmanskonferensen .
Men han gör samma sak själv .
Vi diskuterade och var eniga , utom PPE-gruppen och den liberala gruppen , och jag noterade t.o.m. , det minns ni säkert kära ordförandekolleger , att frågan inte handlar om huruvida ni är för eller emot Todinskatten , utan om ni vågar höra vad kommissionen och rådet tycker om den .
Det är inte för mycket begärt .
Jag upprepar därför förslaget att behålla denna muntliga fråga till kommissionen och rådet för att en gång för alla få veta vilken inställning dessa två instanser har till denna relativt blygsamma begäran , som ändå skulle utgöra en viktig signal till allmänheten , särskilt med tanke på den oro som uppstod efter den misslyckade konferensen i Seattle .
Vi skall rösta om begäran från PPE-DE-gruppen som syftar till att stryka den muntliga frågan om kapitalskatt från föredragningslistan .
( Parlamentet avslog begäran med 164 röster för , 166 emot .
7 ledamöter avstod från att rösta . )
Fru talman !
Jag skulle vilja tacka Poettering för att han just gjort reklam för denna debatt .
Tack .
Fru talman !
Jag undrar om även min röst har räknats , trots att den inte kunde avges på elektronisk väg , eftersom jag inte har något kort ?
Jag röstade " för " .
Om man lägger till de två kolleger som yttrat sig blir resultatet ...
Fru talman !
Ordförandeskapet har redan meddelat resultatet från omröstningen .
Det finns inget utrymme för några ändringar .
( Applåder ) Kära kolleger !
Ännu en gång vill jag påpeka att alla måste ha sitt kort på måndagen .
Det är tydligt att vi har ett problem här .
Jag måste därför fatta ett beslut .
Jag har också glömt mitt kort och jag skulle ha röstat emot .
Jag anser därför att den muntliga frågan kvarstår på föredragningslistan .
( Applåder ) Det är sista gången vi tar hänsyn till att ni glömt korten .
Jag hoppas att alla har förstått och vi skall se till att alla får veta det .
( Applåder ) Ja , den munliga frågan kvarstår på föredragningslistan och , ja , talmannen har rätt att rösta , liksom hon har rätt att också glömma sitt kort .
Vi fortsätter nu med övriga ändringar i föredragningslistan .
Fru talman !
Under den tidigare omröstningen - och jag kommer att följa ert utslag i denna fråga - rörande frågan om kommissionens strategiska plan , sade jag att jag ville uttala mig före omröstningen på min grupps vägnar .
Så blev inte fallet .
Jag skulle uppskatta om jag vid denna punkts avslutande kunde få avge en röstförklaring på min grupps vägnar .
Detta är en viktig fråga .
Det skulle vara användbart för kammarens räkning att upplysa om hur folk uppfattar vad vi just gjort mot bakgrund av deras egen politiska analys .
Fru talman !
Jag skall inte ta upp debatten på nytt , men även jag hade begärt ordet för att ta ställning till herr Barón Crespos begäran .
Ni lät mig aldrig komma till tals .
Det beklagar jag , men omröstningen har genomförts , beslutet har fattats , alltså får det vara .
Jag är ledsen , herr Hänsch och herr Cox , jag såg inte att ni hade begärt ordet .
Jag tror ändå att ståndpunkterna är tydliga och de kommer att bekräftas i protokollet .
När vi i morgon justerar protokollet från dagens sammanträde kan de kolleger , som då anser att ståndpunkterna inte förklarats tillräckligt tydligt , begära ändringar .
Jag tror att det är ett bra sätt .
Naturligtvis kommer man i protokollet från morgondagens sammanträde att ta hänsyn till alla kompletterande förklaringar .
Jag tror att det är bättre än att nu genomföra röstförklaringar som kommer att leda mycket långt .
Vad säger ni om det , herr Cox och herr Hänsch ?
Fru talman !
Om omröstningsregistreringen på ett korrekt sätt visar hur min grupp röstade , skall jag och kan jag inte protestera mot denna .
Om ert utslag innebär att jag inte kan avge en röstförklaring , accepterar jag detta men med reservation .
Vi skall alltså vara mycket noggranna vid upprättandet av protokollet .
Det är vi för övrigt alltid .
Om det inte återger ståndpunkterna tillfredsställande , kan vi eventuellt ändra i det .
( Arbetsplanen fastställdes med dessa ändringar . )
 
Säkerhetsrådgivare för transport av farligt gods Nästa punkt på föredragningslistan är andrahandsbehandlingsrekommendation ( A5-0105 / 1999 ) av Koch , för utskottet för regionalpolitik , transport och turism om rådets gemensamma ståndpunkt inför Europaparlamentets och rådets direktiv om harmoniseringen av examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg eller inre vattenvägar ( C5-0208 / 1999 - 1998 / 0106 ( COD ) ) . .
( DE ) Ärade fru kommissionär , ärade fru talman , kära kolleger !
Jag välkomnar utan förbehåll rådets gemensamma ståndpunkt i strävan mot att skapa en enhetlig utbildning av säkerhetsrådgivare för transport av farligt gods på landsväg , järnväg eller inre vattenvägar .
För det första : vi var tvungna att formellt börja arbeta för att kraven enligt direktiv 96 / 35 / EG skulle uppfyllas , enligt vilka medlemsländerna förpliktigas att vid hantering av farligt gods ta hjälp av ombud resp. säkerhetsrådgivare liksom att organisera utbildning , kurser och examination för dessa personer , utan att utföra detta explicit .
För det andra : genom direktivet uppnår vi a ) bättre säkerhet , såväl under transport som under omlastning av farligt gods ; b ) minskad snedvridning av konkurrensen till följd av de mest skilda nationella utbildningsstrukturer och utbildningskostnader liksom c ) lika villkor för säkerhetsrådgivare på den europeiska arbetsmarknaden .
För det tredje garanterar vi med direktivet såsom det nu föreligger som gemensam ståndpunkt , särskilt i och med att det uteslutande inskränks till miniminormer , en hög grad av flexibilitet och ringa reglering från Europeiska unionens sida , och vi bidrar till stort egenansvar för medlemsländerna .
Allt detta kan vi varmt välkomna i enlighet med subsidiaritetsprincipen .
Jag anser att våra ändringsförslag från första behandlingen har fått vederbörlig uppmärksamhet .
De antogs , andemeningen förverkligades eller också föll de bort på grund av att aktuella europeiska bestämmelser inte infördes , t.ex. ett sanktionssystem mot överträdelser eller en komplicerad blockbildning av frågekomplex .
Jag ber om samtycke till det ena enhälligt godkända ändringsförslaget från utskottet för regionalpolitik och transport , vilket gäller det tidsmässiga införlivandet av direktivet .
I och med att vi inte ger medlemsstaterna något specifikt datum för införlivandet av direktivet utan godkänner en tidsfrist på tre månader från direktivets ikraftträdande , inför vi en flexibilitetsklausul som garanterar ett omedelbart införlivande .
Jag ber om samtycke .
Fru talman !
Vi varken kan eller får finna oss i att allt oftare höra talas om olyckor där stora skador uppstår på våra vägar , men också på järnväg eller inre vattenvägar , inte bara , men också därför att berörda personer inte tar transporten av farligt gods på tillräckligt stort allvar eller därför att okunskap eller bristande utbildning av förarna eller andra ansvariga för de olika kommunikationsmedlen alltför ofta har förvandlat en liten olycka till en stor katastrof .
Jag som österrikare , men jag tror att det gäller oss alla , har fortfarande den katastrof i färskt minne som förra året kostade många människor livet i Tauerntunneln , där det tog många månader av ett enormt ekonomiskt pådrag att bygga upp vad som förstördes vid branden .
Den månadslånga renoveringen skar av denna viktiga trafikled mellan Europas norra och södra delar .
Den omväg för trafiken som detta medförde innebar för många tusen EU-medborgare en påfrestning på gränsen till det uthärdliga .
På sina håll i mitt land var det ett rent helsike .
Förebyggande åtgärder måste bli vårt svar på dylika katastrofer , och med föreliggande direktivförslag skapar vi en viktig grund för att välutbildade säkerhetsrådgivare skall kunna stå till förfogande för att i tid göra det rätta .
Vi får faktiskt inte nöja oss med att skapa en europeisk lag i akt och mening att skapa höjd säkerhet .
Vi måste även konsekvent ge akt på att medlemsstaterna genomför våra riktlinjer inom föreskriven tidsram , och ännu viktigare , vi måste ge akt på att de sedan verkligen tillämpas också .
Inte ännu ett område där vi i efterhand måste beklaga den bristande verkställigheten , tack .
Jag skulle vilja ta upp en sista punkt : Vi får ingalunda nöja oss med att lappa ihop ännu ett hål i säkerhetsnätet och blunda för att det återstår mycket mer att göra på området transportsäkerhet i Europa .
Vidare kräver jag och ber närvarande ansvarig kommissionär att så snart som möjligt lägga fram ett dokument som sörjer för bättre säkerhet i framtida tunneltrafik så att vi slipper uppleva fler katastrofer av denna vidd här i Europa !
Fru talman !
Låt mig först och främst tacka Koch för hans betänkande , i vilket han på ett mycket seriöst sätt behandlat frågan om transportsäkerhet .
Han behandlar frågan om harmonisering av examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg och inre vattenvägar .
Jag gratulerar honom till hans utmärkta betänkande .
Transportsäkerheten har tråkigt nog diskuterats i nyheterna nyligen : Tågkraschen vid Paddington i London , den fruktansvärda tågkraschen i Norge , de två flygkrascherna där EU-medborgare fanns ombord och naturkatastrofen utanför Bretagnes kust efter Erikas haveri - som alla skett inom de senaste fyra månaderna - påminner oss om att transportsäkerheten aldrig kan tas för given och de som ansvarar för att skydda allmänheten måste vara mycket motiverade och mycket kvalificerade .
Föredraganden har påpekat för kammaren att rådet i sin gemensamma ståndpunkt har godkänt sex av parlamentets tio ändringsförslag som lades fram vid första behandlingen , och att andemeningen i parlamentets övriga ändringsförslag har behållits .
Min grupp vill därför stödja den gemensamma ståndpunkten och ser fram emot antagandet av lagstiftningen , vilken kommer att ge oss ytterligare ett instrument i vår kamp för att göra transporterna i Europeiska unionen så säkra som möjligt .
När det gäller säkerhet kommer min grupp alltid att stödja initiativ som avser att förbättra transportsäkerheten .
Som händelserna under den senaste tiden visat , har vi fortfarande mycket arbete kvar på detta område .
Fru talman !
I detta parlament uppmärksammas regelbundet , med rätta , hur viktig transportsäkerheten är .
De alltjämt ökande mängder gods som transporteras genom Europa medför medvetet och omedvetet allehanda risker för personalen och samhällsomgivningen .
De som måste hantera dessa risker måste därför uppfylla höga krav .
De normer för detta som fastlagts i ett annat direktiv , 95 / 35 / EG , förefaller vara tillräckligt adekvata för att på ett ansvarigt sätt ge råd om hur transporter av farligt gods skall organiseras .
Det gläder mig att vi också nått samförstånd med rådet i fråga om minimikraven för deras examen , även om jag hellre hade sett att enhetliga fasta normer kommit till stånd , så att examensbevisen är lika internationellt sett .
Men det har visat sig att detta inte går att uppnå .
Slutligen , ändringsförslaget som föredraganden föreslår är inte mer än logiskt , och därför kan jag också helhjärtat stödja detta .
Herr talman , fru kommissionär , ärade kolleger !
Först vill jag gratulera min kollega Koch till hans betänkanden , som måhända är tekniska rapporter , men som har mycket stor betydelse för säkerheten .
Jag vill endast göra några små anmärkningar .
Först vill jag be fru kommissionären - och jag är övertygad om att min önskan faller i god jord - att ägna säkerhetsfrågan större uppmärksamhet , vare sig det gäller på vägar , på inre vattenvägar eller på havet .
När jag inser att den första begäran gjordes till kommissionen den 19 mars 1998 och att vi behandlar frågan här i dag - trots att parlamentet reagerade relativt snart - då tycker jag att tidsrymden är något för lång .
Nu är detta inte enbart kommissionens fel , men jag tycker att vi måste reagera snabbare för att få till stånd en standardisering även här .
Den andra punkten nämndes just : minimireglerna .
Jag är principiellt av den åsikten att vi på många transportområden borde eftersträva ökad flexibilitet samt regelverk som gäller land för land .
När det gäller säkerheten är jag dock något skeptisk , eftersom säkerheten i låt oss säga Sverige i princip inte skiljer sig från säkerheten i Tyskland , Italien eller Österrike .
Jag kan leva med dessa minimiregler , men jag ber kommissionen att verkligen uppmärksamt följa händelseutvecklingen .
Om den här typen av flexibilitet i vissa länder skulle leda till bristfälliga bestämmelser , då bör vi genomföra ytterligare standardiseringar .
Den tredje punkten har även den nämnts .
Jag kommer ju , precis som min kollega Rack , från ett transitland , där denna fråga spelar en särskild roll .
Vi skall inte försämra konkurrensvillkoren ensidigt för vissa länder och förbättra dem för länder som Österrike eller andra transitländer .
Men jag anser att vi bör göra allt för att hålla transporten av farligt gods på så låg nivå som möjligt , och det i alla länder , transitland eller inte .
Herr talman !
Jag vill börja med att gratulera föredragande Koch till hans utmärkta arbete och hans konstruktiva samarbete med kommissionen när det gällt att förbättra texten , föredra detta betänkande och förslag ; slutligen finns det endast ett ändringsförslag beträffande examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg eller inre vattenvägar .
Vi anser att samarbetet är av stor betydelse , de gemensamma insatserna från de båda institutionerna - parlamentet och kommissionen - och samarbetet med utskottet för regionalpolitik , transport och turism , med transportgruppen närmare bestämt , fungerar alldeles utmärkt .
Den gemensamma ståndpunkten inbegriper praktiskt taget alla ändringsförslag som har godkänts av kommissionen , examineringskraven för säkerhetsrådgivare har harmoniserats och , i andra behandlingen , kan vi godkänna ändringsförslaget med ett datum som är mer realistiskt än det datum som kommissionen föreslog i början , med tanke på att vi redan har debatterat den här frågan i många år .
Jag vill också kort tacka de olika parlamentsledamöterna för deras insats och tala om för er , mina damer och herrar , att kommissionen prioriterar säkerheten på transportområdet .
Och Simpson har alldeles rätt i det han sade , att man aldrig får betrakta processen som slutförd , som avklarad eller som färdig .
Processen med ett utökande av marginalerna , av säkerhetsgarantierna vid transport är en process som måste förbättras dag för dag .
I den bemärkelsen vill jag också kort ta upp problematiken med tunnlarna , som Rack och Swoboda hänvisade till , och som utan tvekan är en mycket känslig fråga för Österrikes del , och vi måste därför bemöda oss om att förbättra säkerheten .
Vid en av de större olyckor som inträffat på senare tid , var inte det transporterade godset farligt i sig .
Margarin och några kilo målarfärg , som i princip inte utgjorde någon risk , kom att orsaka en riktig katastrof .
Därför måste man fundera över hur man ytterligare kan skärpa de krav som garanterar en maximal säkerhet .
Avslutningsvis vill jag säga att säkerheten måste iakttas vid alla typer av transporter .
Den här veckan skall vi hålla en debatt där vi talar om säkerheten vid sjötransporter , till följd av katastrofen med Erika , och vi kommer under det här året att få diskutera målsättningen i fråga om säkerhet vid flygtransporter .
Mina damer och herrar , jag vill påpeka att säkerheten är ett mål som prioriteras av kommissionen .
Och som jag kommer att säga i debatten om Erika , får vi inte vänta tills det inträffar en katastrof innan vi tar itu med säkerhetsaspekten .
Låt oss i stället ta oss an frågan utanför sådana situationer som inte utgör annat än ett bevis på hur brådskande det är med en effektiv lösning på denna typ av problem .
Jag vill än en gång rikta ett tack till alla som har medverkat och då i synnerhet föredragande Koch .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Transport av farligt gods på väg Nästa punkt på föredragningslistan är betänkande ( A5-0104 / 1999 ) av Koch för utskottet för regionalpolitik , transport och turism om Europaparlamentets och rådets direktiv om ändring av direktiv 94 / 55 / EG om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg [ KOM ( 1999 ) 158 - C5-0004 / 1999 - 1999 / 0083 ( COD ) ] . )
Herr talman , ärade fru kommissionär , kära kolleger !
Det direktiv som trädde i kraft den 1 januari 1997 om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg innehåller en del övergångsbestämmelser , vars giltighet är temporär och knuten till att CEN , alltså Europeiska standardiseringskommittén , utarbetar bestämda regler .
De dröjsmål som har uppstått i CEN : s arbete leder nu till problem med införlivandet av direktivet .
Framför allt kan bilagorna inte anpassas i takt med den tekniska och industriella utvecklingen .
Jag beklagar detta , för nu måste vi göra det arbete andra inte har gjort .
I så måtto accepterar jag föreliggande förslag om ändring av direktiv 94 / 55 / EG , vilket skall diskuteras i dag .
Om Europeiska unionen avstår från att gripa in skulle detta tvinga medlemsstaterna att ändra sina inhemska rättsliga bestämmelser för en kort period , nämligen tills CEN : s arbete har slutförts , vilket drar med sig onödiga kostnader och förvirring .
Den ändring av direktivet som i dag står på föredragningslistan innebär alltså ingen förändring i den standardisering av transport av farligt gods som gemenskapen har i dag .
Genom denna utvidgas däremot övergångsbestämmelserna genom att gällande datum skjuts upp , de bestämmelser som inte längre är relevanta stryks och den innebär att förfarandet regleras vid a ) ad hoc-transporter av farligt gods liksom b ) införandet av mindre stränga nationella bestämmelser , särskilt vad gäller transport av mycket ringa mängder farligt gods på geografiskt sett mycket strängt avgränsade områden .
Därmed ligger ändringen av direktivet helt i linje med subsidiaritetsprincipen : medlemsländerna får större befogenheter .
EU-kommissionen avgör huruvida medlemsländerna kan införa egna särskilda bestämmelser .
Kommissionen stöds efter regleringsförfarandet av ett expertutskott för transport av farligt gods .
Detaljerna för hur dessa befogenheter som anförtrotts kommissionen skall utövas har ändrats i rådets beslut från juni 1999 .
Det förslag till ändring av direktivet gällande transport av farligt gods på väg , som skall diskuteras i dag , är dock från maj 1999 och har därför ännu inte kunnat ta hänsyn till det aktuella kommittéförfarandet .
De framlagda och av utskottet enhälligt godkända ändringsförslagen åberopar i två fall just detta förändrade kommittéförfarandet .
Vi skulle vilja säkerställa att det redan i motiveringen hänvisas till detta och att den icke entydigt formulerade tidsfristen , inom vilken rådet måste fatta beslut , fastställts till högst tre månader .
Därutöver hänvisas det till nödvändigheten av ökad öppenhet .
Ett annat ändringsförslag tillåter medlemsländerna att införa skärpta krav , framför allt för vakuumtankar , för arbete resp. transport vid temperaturer på under minus 20 º C. Detta är särskilt intressant för de nordeuropeiska regionerna .
Ett sista ändringsförslag skall göra det tillåtet att fortsätta använda de tankar och tankfordon som tagits i bruk mellan den 1 januari 1997 och ikraftträdandet av detta direktiv , under förutsättning att de konstruerats och servats på vederbörligt sätt .
Även om jag är medveten om att detta endast är ett litet steg mot ökad transportsäkerhet ber jag er anta betänkandet .
Herr talman , bästa kolleger !
Gott nytt år och gott nytt millennium !
Det är första gången jag talar vid plenarsammanträdet och detta är spännande , i viss mån likt den första kärleken , men den första kärleken varade dock längre än två minuter .
Jag skulle kort vilja kommentera kommissionens förslag till ändring av direktivet om transport av farligt gods på väg .
Det är bra att detta direktiv utfärdas nu eftersom medlemsstaterna i annat fall skulle tvingas att ändra sina nationella bestämmelser för en mycket kort tid , en övergångsperiod , vilket i sin tur bara skulle förorsaka onödiga kostnader och än en gång öka allmänhetens grämelse över EU : s byråkrati .
I kommissionens förslag har man emellertid inte tagit hänsyn till alla aspekter , som till exempel de nordliga regionernas kalla klimat .
Därför har jag föreslagit några ändringar , som godkänts i vårt utskott , till kollegan Kochs i och för sig utmärkta betänkande .
Mina ändringsförslag gäller köldbeständigheten hos de tankar som används för transport av dessa farliga ämnen .
Enligt kommissionens förslag skulle det räcka med minus tjugo grader ; vid Medelhavet har man svårt att föreställa sig att temperaturen i Lappland skulle kunna sjunka betydligt lägre .
Även i Lappland stödjer man EU , låt oss därför även komma ihåg dem som bor där .
Således föreslår jag att köldgränsen skall sänkas till minus fyrtio grader .
Detta är också nödvändigt för att bibehålla nuvarande säkerhetsnivå i de nordliga områdena .
Jag hoppas att mina förslag beaktas vid omröstningen i morgon .
Herr talman !
Tillåter ni att jag först av allt uttrycker min respekt för ert sätt att klara det flygande bytet på ordförandebänken under debatten för en stund sedan .
Det var lysande .
Till saken : Jag anser att Europas medborgare måste kunna lita på att det som transporteras på Europas vägar , järnvägsnät osv . , även om det är farligt gods , transporteras så säkert som möjligt .
Direktivet är ett bidrag till detta .
Vad vi gör här i dag är i grund och botten ett irritationsmoment .
Föredraganden Koch , som vi tackar för det arbete han har utfört , har påpekat att i princip allt redan hade kunnat komma längre om det inte hade varit för försummelsen från CEN , som är mycket senfärdig med att upprätta och anpassa riktlinjen .
Därför kan vi bara hoppas - och denna vecka helst besluta om - att vi år 2001 äntligen får en gemensam reglering av transporten av farligt gods på väg , så att vi får en gnutta rättssäkerhet här inne och en gnutta ökad säkerhet där ute på våra vägar .
Fru kommissionär , herr talman !
Låt mig börja med att tacka herr Koch för hans betänkande , som är utmärkt , och jag har heller inte alltför mycket att tillägga .
Jag vill dock ta tillfället i akt och påpeka att det inte bara är i Indien , som jag just återvänder ifrån , utan också i EU som risktransporter fortfarande medför stora problem .
Vi behöver bara tänka på den svåra olyckan i Mont Blanc-tunneln för runt ett år sedan - även Tauerntunneln hör dit .
Vi ser att det alltid är i områden där själva naturen skapar svårigheter - dimma , stormar , kyla - och framför allt i de trånga passen i alperna som det i sammanhanget fortfarande kan uppstå stora problem .
Jag pläderar generellt för att farligt gods i större utsträckning skall flyttas över till järnvägen .
I förebyggande syfte måste rätt lösning för framtiden finnas med redan i planeringen av framtida sträckor - järnväg eller också motorväg .
Tänk bara på Brenner-Basistunneln som ännu inte har diskuterats på djupet .
Jag vill också understryka att transportproblematiken är en av nyckelfrågorna inom EU och be kommissionen ta detta på allvar .
För att förbättra funktionaliteten måste vi föra mycket mer intensiva och återkommande diskussioner om hur transporter kan undvikas , om tung trafik till järnväg , om vägavgifter och privatisering av järnvägen .
När jag tänker på att utvidgningen österut kommer att föra ytterligare några problem med sig så inser vi alla att EU : s trovärdighet i framtiden även kommer att bero på om och hur vi lyckas reglera trafiken .
Herr talman !
Det betänkande som vi här behandlar innebär i sig inga stora förändringar .
De flesta av ändringsförslagen är av enbart teknisk natur .
Det är dock värt att understryka att varje gång som vi fattar denna typ av beslut är det bra ur ett brett miljöperspektiv , och det är bra därför att det skapar bättre förutsättningar för den inre marknadens möjligheter att fungera .
Det transporteras runtom i EU mycket stora mängder farligt gods både på vägar , järnvägar och på haven .
Det gör att det är nödvändigt med ordentliga regler för hur detta skall fungera .
På område efter område får vi nu gemensamma minimiregler för medlemsländerna .
Det är utomordentligt positivt , och det finns anledning att tacka föredraganden , Koch , för det arbete som han har lagt ned på detta ärende .
Detta är också viktigt när det gäller förutsättningarna för den inre marknaden .
Om vi skall få en gemensam transportmarknad att verkligen fungera , är det viktigt , inte bara att vi har regler , utan också att dessa regler så långt som möjligt är gemensamma .
Jag vill avslutningsvis gärna kommentera en tredje sak som också är väsentlig , nämligen ett ändringsförslag framlagt av ledamoten Ari Vatanen .
På många sätt skiljer sig förutsättningarna från ett medlemsland till ett annat .
Genom att godkänna detta ändringsförslag , tar vi hänsyn till att det i de norra delarna av unionen kan vara mycket kallt .
Det gör att det är nödvändigt att också ta hänsyn till hur material och förpackningar påverkas av en sådan kyla .
Herr talman , det är positivt att vi i denna reglering också kan vara flexibla .
Det är min förhoppning att kommissionen kan acceptera denna ändring .
Herr talman !
Jag vill tacka inte bara kollegan Koch , utan också vice ordföranden i kommissionen för hennes klara och entydiga ställningstagande för säkerheten på transportområdet och prioriteringen av säkerheten .
Koch har producerat ett bra betänkande , emedan det inte har kommit ut mycket av arbetet på CEN eller inom ramen för Förenta nationernas ekonomiska kommission för Europa .
Jag vill fråga vice ordföranden om hon i dag kan säga oss hur läget är när det gäller standardiseringssträvandena i dessa båda organisationer samt om EU har möjlighet att snabba på standardiseringssträvandena enligt enklast möjliga principer .
För det står klart att även om vi inför fantastiska bestämmelser här inom Europeiska unionen så gör trafiken inte halt vid dessa gränser , den överskrider dem .
Därför är det säkerligen meningsfullt med mer långtgående , nämligen regionalt sett mer långtgående regleringar .
Om det inte är möjligt att svara på detta i dag , vore det då möjligt att utskottet får ett skriftligt meddelande om hur läget ser ut och hur det står till med förhandlingarna mellan CEN och FN : s ekonomiska kommission för Europa ?
Herr talman !
Jag upprepar mina gratulationer till herr Koch för hans arbete med det här betänkandet , som på sätt och vis har blivit ett komplement till den debatt vi höll i oktober månad om transport per järnväg .
Alla beklagar vi att Europeiska standardiseringskommittén ( CEN ) inte har haft förmåga att inom de uppställda tidsramarna slutföra den ändring av de bestämmelser som krävs för en lämplig harmonisering inom Europeiska unionen .
Den här debatten och ändringen av det nu gällande direktivet gör att vi kan ta med andra fakta som visar på mångfalden i vårt Europa .
För en stund sedan talade Vatanen om låga temperaturer , inte bara om 20 minusgrader utan om 40 minusgrader .
Naturligtvis godkänner vi det ändringsförslaget , han har helt rätt , och jag anser att man bör ta med konkreta omständigheter som visar på det varierade klimatet i Europeiska unionen , som i vissa fall omvandlas till specificeranden och konkreta krav när man tittar på standardiseringar och karakteriseringar av teknisk art .
Vad beträffar Swobodas uttalanden om CEN : s verksamhet , kan jag tala om att vi har uppmanat dem att påskynda arbetet så mycket som möjligt , för det skulle vara illa om vi , trots den nya fristen , skulle stå inför samma problem om drygt ett år på grund av att arbetet inte har slutförts .
Slutligen , herr talman , kan sägas att vi har lyft fram de grundläggande problem som rättfärdigar en ändring av direktivet , vi har talat om förseningen från CEN : s sida , om ändringar av vissa bestämmelser , om sambandet mellan direktivets text och innehållet i bilagorna , om behovet av en närmare precisering .
Alla bidrag från parlamentets utskott och föredraganden Koch , som har omvandlats till olika ändringsförslag , närmare bestämt i fyra , har antagits av kommissionen .
Vi godkänner således de fyra ändringsförslag som har lagts fram för oss .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Samordning strukturfonderna / sammanhållningsfonden Nästa punkt på föredragningslistan är betänkande ( A5-0108 / 1999 ) av Schroedter för utskottet för regionalpolitik , transport och turism om meddelandet från kommissionen om samordning av strukturfonderna och Sammanhållningsfonden - Riktlinjer för programmen för perioden 2000-2006 [ KOM ( 1999 ) 344 - C5-0122 / 1999 - 1999 / 2127 ( COS ) ] . .
( DE ) Herr talman , fru kommissionär !
Ah , herr kommissionären är här , och jag som trodde att ni inte skulle komma .
Välkommen till parlamentet !
Kära kolleger !
Vi kan inte blunda för att vinsterna på den europeiska hemmamarknaden är koncentrerade till de rika regionerna och inte ens där kommer alla delar av befolkningen till godo .
Hur länge skall vi egentligen acceptera en utveckling som resulterar i ökade klyftor mellan fattiga och rika regioner ?
Medan det i den femte rapporten om situationen i regionerna meddelas att arbetslösheten i de fattiga regionerna var sju gånger så hög som i de rika regionerna , talas redan i den sjätte rapporten om en åtta gånger så hög arbetslöshet , trots att anslag från de europeiska strukturfonderna flyter in i regionerna .
Därför blir naturligtvis ingen förvånad över att det redan i inledningsskedet av den nya strukturfondförordningen reses krav på att resurserna skall användas på ett mer effektivt och koncentrerat sätt i den europeiska målsättningen att nå hög sysselsättningsnivå och bestående utveckling , för att endast nämna några .
Parlamentet , men framför allt medlemsstaterna ställde massiva krav på förbättringar .
Detta föll emellertid relativt snart i glömska i och med att kommissionen utvecklade det nya instrumentet för detta - riktlinjerna - och ville göra kraven på effektivitet , koncentration och enklare förvaltningsförfaranden mer bindande vid tillämpningen av de europeiska strukturfonderna .
Då åberopade medlemsländernas regeringar subsidiaritetsprincipen och ville helt enkelt få sig pengarna tillskickade .
Av toppmötet i Berlin 1999 blev sålunda endast riktlinjernas vägledande karaktär kvar .
Men dessa förpliktar åtminstone kommissionen att endast godkänna program som leder till att de europeiska målen faktiskt kan uppnås .
Även om jag tvivlar på att detta vägledande instrument verkligen räcker till för att uppnå effektivitet och koncentration och för att i realiteten förverkliga de europeiska målen , så kvarstår det faktum att riktlinjerna kommer att spela en central roll i förhandlingarna om gemenskapsstödramen .
Och det måste de göra om man på europeisk nivå vill bli tagen på allvar !
Parlamentet hade ingen möjlighet att gå in på innehållet i riktlinjerna , eftersom man rådfrågades först när mandatperioden redan var över .
Nu när programplaneringsfasen är så långt framskriden är det knappast meningsfullt att ta tillbaka alltihop .
Därför koncentrerar jag mig , med utskottets goda minne , i mitt betänkande på instrumentets strategiska karaktär .
För det första : i betänkandet granskas resultatet av instrumentet i sig .
För det andra : det avslöjar bristerna i kommissionsdokumentet .
Så har till exempel partnerskapet rätt och slätt glömts bort i den centrala delen av strukturfonderna .
Förgäves letar man i dokumentet efter den centrala princip som uppmanar medlemsstaterna att på hemmaplan arbeta fram program tillsammans med kommunerna och regionerna men också med de lokala aktörerna , ekonomiska och sociala organisationer , icke-statliga organisationer , fackföreningar , företagarföreningar , kvinnoförbund , aktionsgrupper , sysselsättningsinitiativ .
Frågan varför detta glömdes bort har den dag som i dag är ännu inte besvarats .
Här ställer parlamentet centrala krav .
Parlamentet förväntar sig att kommissionen endast bifaller program som har arbetats fram i ett sådant partnerskap .
Jag är förvånad , kära kolleger från den konservativa gruppen , att jag så plötsligt över en natt finner ändringsförslag enligt vilka man vill stryka de decentralistiska ansatserna .
Jag kan bara säga , ta med förslagen till era regioner och förklara för era väljare varför den europeiska principen om decentralisering inte skall förverkligas ute i regionerna .
Jag lovar att ni inte kommer tillbaka helskinnade .
Det får inte gå till så att vi sitter här och utarbetar principer , men när det gäller genomförandet så gör var och en vad hon eller han vill .
En kommentar i förbifarten till regeringen i mitt land där man helt enkelt vill ignorera den horisontella gemenskapspolitiken när det gäller miljöskydd och inte tyckte sig behöva följa direktivet om bevarande av livsmiljöer samt vilda djur och växter : jag uppskattar att kommissionen är hård på den punkten .
Och därmed är jag inne på den sista punkten .
Riktlinjerna måste bli en konkret måttstock för huruvida artikel 1 i förordningen efterlevs eller inte .
Jag förväntar mig att kommissionen kommer att se till att riktlinjerna , som faktiskt erbjuder tillräcklig flexibilitet , verkligen får utgöra själva måttstocken för förhandlingarna .
Vi företräder den europeiska ståndpunkten .
Det innebär att lika stor hänsyn måste tas till beständigheten i transportpolitiken som till andelen kvinnor i produktionen liksom till det faktum att varje program föreskriver omfattande bidrag , vilket möjliggör en bestående utveckling i städerna och pilotprojekt för landsbygdsområdena .
Jag förväntar mig att detta får bli resultatet av gemenskapsstödramen och att ni inte säckar ihop igen .
För hur skall vi annars få arbetslöshetssiffrorna att sjunka om vi avvaktar igen , om vi återigen försöker fuska oss dit ?
Vi kan inte avvakta !
Det här är de sista åren som vi har möjlighet att driva den europeiska strukturpolitiken med så omfattande finansiering .
Därefter tillkommer många nya länder , och då blir vi hur som helst tvungna att skapa bättre , mer effektiva och koncentrerade strukturer .
Och det är bara början .
Det är därför jag förväntar mig att kommissionen i förhandlingarna skall ta parlamentets krav på allvar och verkligen omsätta den europeiska ståndpunkten i handling och därmed äntligen ge en progressiv regionalpolitik chansen .
Herr talman !
Det är särskilt tillfredsställande för mig att hålla mitt första tal i Europaparlamentet om vad som anses vara den viktigaste frågan i den del av Förenade kungariket som jag företräder i detta parlament , dvs .
Wales .
Huvuddelen av Wales har , som ni känner till , erkänts mål 1-status enligt strukturfondsprogrammen .
Det är helt klart så att många i Wales förlitar sig på Europeiska unionens strukturfondsprogram när det gäller att lindra en del av de enorma svårigheter som vi utan tvekan står inför .
Vi har sett att fattigdomen ökar i Wales ; och har ökat ytterligare sedan 1997 .
Vi har sett klyftan mellan rika och fattiga vidgas .
Vi förlitar oss därför på strukturfondsprogrammen , inte bara för att få till stånd en industriell omstrukturering , utan också för att få till stånd en bredare förbättring av hela den ekonomiska basen i Wales .
Vad som emellertid är djupt skadligt för oss , är tron att beviljandet av medel från strukturfonderna är något som , på sätt och vis , varit en framgång för regeringen .
Det är tråkigt nog bara ett erkännande av de mycket stora svårigheter som Wales står inför .
Detta är skälet till varför jag vill betona vissa av de frågor som jag anser att kommissionen måste prioritera .
Vi vänder oss till kommissionen för att ta itu med frågor som har att göra med kompletterande medel .
Vi är missnöjda med det faktum att dessa siffror på något sätt verkar har gömts i Förenade kungarikets siffror .
Vi vänder oss också till kommissionen för att se till att det finns matchande finansiering för projekten .
Vi vänder oss till den för att utmana den brittiska regeringen , för att se till att privata sektorn - som antagligen måste stå för den största delen av utgifterna inom strukturfonderna - deltar vid planeringsstadiet .
Vi uppmanar , till sist , kommissionen att se till att pengar från strukturfonderna används på ett öppet och väl redovisat sätt .
Alltför mycket av vad som sker i detta parlament är inte öppet och väl redovisat .
Detta är ett område inom vilket kommissionen kan hjälpa Wales på ett avgörande sätt .
Herr talman !
Vårt utskott studerar dessa frågor ur många olika synvinklar , men först skall jag tala om forskningens synvinkel .
Vi ser mycket positivt på att föredraganden i sina egna slutsatser inkluderat vårt utskotts förslag om att man borde utvidga forskningsinfrastrukturen i sammanhållningsländerna genom att placera ut högskolor och läroanstalter så att de bättre tjänar invånarna i mindre utvecklade regioner och gör det lättare för utbildade personer att stanna kvar i sin hembygd .
Detta kan ske genom myndighetsåtgärder , och en sådan decentralisering av den högre utbildningen är utan tvivel nyttig för att utjämna utvecklingen .
En annan fråga som vi uttryckligen skulle vilja belysa ur en industripolitisk synvinkel är att vi gärna sett att kommissionen fäst större uppmärksamhet vid effekterna av ökad användning av tjänster , elektronisk handel och Internet när den planerade samordningen av strukturfonderna och Sammanhållningsfonden .
Tidigare fanns det ett större samband mellan fattigdom / rikedom och näringsstrukturen .
Rika var de områden där det fanns arbetstillfällen inom industrin , men i dag har dessa områden kanske blivit till en belastning och kan vara fattiga , vilket gör att man också måste satsa på nya verksamhetsgrenar , på så kallad elektronisk produktion och tjänsteproduktion , eftersom detta är framtidens verksamhetsgrenar .
Det ansvariga utskottet har enligt min mening inte i tillräcklig utsträckning tagit hänsyn till detta i sitt betänkande , varför jag å utskottets för industrifrågor vägnar önskar rikta kommissionens uppmärksamhet på denna fråga .
Till slut skulle vi i egenskap av utskott för energi ha önskat att man i ännu högre grad framhållit stödet för förnybara energikällor från Sammanhållningsfonden och regionala utvecklingsfonden , och därigenom hade man med hjälp av samordning kunnat öka användningen av förnybara energikällor så att energiprogrammets otillräckliga finansiering kompenserats med dessa mer omfattande penningresurser . .
( EN ) Herr talman !
Jag vill verkligen tacka fru Schroedter för det arbete hon lagt ned i detta sammanhang och förklara för mina kolleger att uttalar mig på min kollega Flautres vägnar , som följde detta för utskottet för sysselsättning och socialfrågor , men som tyvärr blivit sjuk .
Jag vill rikta uppmärksamheten på ändringsförslag 1 och 2 , vilka röstades igenom av utskottet för sysselsättning och socialfrågor , men inte godtogs av utskottet för regionalpolitik , transport och turism .
Dessa ändringsförslag behandlar den sociala ekonomin och behovet av att tillhandahålla socialt riskkapital och finansiellt stödja lokala program för utveckling av sysselsättningsmöjligheter och stärkande av den sociala sammanhållningen .
Under årens lopp har parlamentet sett den sociala ekonomin som en viktig och möjlig skapare av arbetstillfällen .
Dessa ändringsförslag överensstämmer också med parlamentets syn att social utslagning är en viktig fråga som kräver konstruktiva åtgärder .
Vi hoppas att de som överväger att förkasta dessa ändringsförslag har mycket kraftfulla skäl att erbjuda både parlamentet och de medborgare som letar efter arbete .
I sitt betänkande pekade också Flautre på ett område inom vilket det i högsta grad saknas samordning , fast detta sannerligen behövs .
I kommissionens förslag hänvisar man till sysselsättningsstrategins fyra pelare och Europeiska socialfondens fem åtgärdsområden .
Men det är särskilt beklagligt att det här saknas specifika riktlinjer , då idén med att sammanlänka hjälp från socialfonden till sysselsättningsstrategin kommer att träda i kraft för första gången under programperioden 2000-2006 .
Man kan säga att denna försummelse ger intrycket att också kommissionen inte har någon idé om hur den skall skapa högsta möjliga samordning mellan hjälp från socialfonden , vilken skall granskas efter tre och ett halvt år , och medlemsstaternas årliga nationella sysselsättningsplaner .
Vi hoppas att kommissionen kan ge oss lugnande besked om att detta var ett förbiseende som man nu skall ta itu med på ett konstruktivt sätt .
Herr talman , herr kommissionär , ärade parlamentsledamöter !
Det förslag som kommissionen har lagt fram av , och därmed uppfyller sitt mandat , betraktar utskottet för jordbruk och landsbygdens utveckling som en vettig utgångspunkt .
Men jag vill här poängtera att denna utgångspunkt visar vilka utmaningar vi nu står inför : att förmå befolkningen att stanna kvar på landsbygden , med de förändringar som håller på att ske inom all ekonomisk verksamhet på grund av jordbrukssektorns allt minskande betydelse som inkomstkälla på landsbygden .
Detta , tillsammans med bristerna i infrastrukturnätet och samhällsservicen , och arbetstillfällena som i regel är få , ofta säsongsbetonade och tämligen likriktade , ökar flykten från landsbygden .
Följderna låter inte vänta på sig .
Det är ungdomarna som försvinner , som utbildar sig och får arbete i städerna , något som påverkar landsbygden på ett negativt sätt .
Denna bristande infrastruktur är också ett hinder för utbredningen av företag och skapandet av nya arbetstillfällen .
Man bör komma ihåg att landsbygden utgör nästan fyra femtedelar av Europeiska unionens yta .
Inom jordbruket finns endast 5,5 procent av alla arbetstillfällen i unionen .
Dessutom driver tre fjärdedelar av alla jordbrukare jordbruk som en deltidssysselsättning och är beroende av ett effektivt tillägg till sina inkomster .
Ett av de främsta och viktigaste målen som vi bör fastställa i Europeiska unionen är därför att bemöda oss om att skapa nya arbetstillfällen på landsbygden , utanför jordbrukssektorn , inom sektorer som landsbygdsturism , sport , kultur , återerövrande av fädernearvet , omvandling av företag , nya tekniker , tjänstesektorn , etc .
Även om jordbruket inte längre har en exklusiv roll fortsätter det att vara viktigt , inte bara för att undvika att landsbygden hamnar utanför i ekonomiskt och socialt avseende och att nya spökstäder uppkommer , utan även för att jordbrukarna har en viktig roll i förvaltningen av territoriet , bevarandet av den biologiska mångfalden och skyddet av miljön .
Därför förespråkar vi att man fastslår en politik för jordbruket och landsbygdens utveckling som överensstämmer med de mål som vi har satt upp och att landsbygden , i början av 2000-talet , skall vara konkurrenskraftig och mångfunktionell , såväl ur jordbrukssynpunkt som beträffande en öppen attityd gentemot olika verksamheter utanför jordbruket .
Det är viktigt att prioritera de allmänna kriterierna för en översiktsplan och befolkningsspridning , och beakta slutsatserna från utskottet för jordbruk och landsbygdens utveckling i fem viktiga avseenden , som endast i viss utsträckning har anammats av utskottet för regionalpolitik , transport och turism under punkterna 16 och 17 .
Slutligen vill jag be kommissionen att dessa fem punkter beaktas vid fastställandet av slutsatserna för de fyra pelarna , för jag anser att bevarandet av befolkningen på landsbygden bör vara ett av Europeiska unionens främsta mål .
Herr talman , herr kommissionär , ärade kolleger !
Jag vill börja mitt anförande med att tacka föredragande Schroedter för hennes insats .
Jag anser att det är ett väl genomarbetat betänkande .
Dessutom vill jag tacka henne för hennes vilja till dialog med de övriga politiska grupperna när det var dags att uppnå en avtalslösning inför denna våg av ändringsförslag , som kanske var fler än man hade räknat med , men dessa speglar i själva verket vikten av det betänkande som vi nu diskuterar .
För oss är det viktigt att de slutsatser som antas av parlamentet beaktas av kommissionen , åtminstone andemeningen av dessa , för annars kan det i den här situation verka som att det vi ägnar oss åt är meningslöst och endast en övning i retorik .
Faktum är att vi anser , och det framgår av ordalydelsen i slutsatserna , att kommissionen bör ta hänsyn till det som beslutas här i parlamentet , i första hand om granskningen av dessa riktlinjer när halva tiden har gått .
I våra ändringsförslag har vi fastslagit hur viktigt det är att man skapar den nödvändiga samordningen mellan strukturfonderna , Sammanhållningsfonden och gemenskapsinitiativen , så att tillämpandet av dessa på bästa sätt , på det mest lönsamma sättet speglar sig i ett successivt utplånande av olikheterna mellan regionerna och i skapandet av sysselsättning , utan tvekan de två viktigaste målsättningarna för de fonder vi talar om .
Och som ett sätt att ge en snabb och effektiv impuls till att uppnå dessa målsättningar , anser vi att det är viktigt att de som skapar sysselsättning medverkar i detta initiativ , de som verkligen är driftiga och de som verkligen kan garantera nya arbetstillfällen , det vill säga företagarna .
Utdelningen av dessa fonder måste i synnerhet komma de mindre och mellanstora företagen till godo .
Om det inte skulle vara fallet , om företagarna känner sig utstötta , om inte företagarna får ta del , och då menar jag inte bara i förvaltningen , utan även i mottagandet av dessa fondmedel , då har vi missat en möjlighet att uppnå våra mål på snabbast tänkbara sätt .
Dessutom är det viktigt att vi för att uppnå dessa , för att övervinna olikheterna mellan regionerna och finna källor till sysselsättning , satsar rejält på de nya teknikerna , på näten för transport och kommunikation och på förnybara energikällor .
Och detta - jag upprepar - med medverkan av de privata företagen som genom att förena sina insatser med insatserna från den offentliga förvaltningen , som ett komplement till denna utan att det ena för den skull skall hindra eller utesluta det andra , är de som kommer att skapa ett rikt samhälle och nya arbetstillfällen .
Herr talman !
Det åligger mig att påminna min kollega , Evans , om varför Wales egentligen erhöll mål 1-status .
Det berodde på den skamliga politik som hans eget parti , de konservativa , förde .
Låt mig också påminna honom om att när hans partiledare , Hague , var Wales utrikesminister , bröt han mot varenda regel rörande kompletterande medel , vilket resulterade i ett skarpt formulerat brev från kommissionsledamot Wulf-Mathies angående föreskrifterna .
Jag kan försäkra er om att den brittiska regeringen känner till sina föreskrifter rörande kompletterande medel för mål 1 .
Jag föreslår att Evans läser bestämmelserna .
Min grupp har lagt fram omfattande ändringsförslag till båda de betänkanden som debatteras i dag .
Jag vill att vi koncentrerar oss på riktlinjernas avgörande roll .
Målet är att tillhandahålla en ram - ett instrument - för stöd och förstärkning av den ekonomiska förnyelsen , för att på ett effektivt sätt använda resurserna i de mest långtgående partnerskapen och att få dessa regioner på rätt köl , så att de kan återhämta sig och få en hållbar utveckling och slutligen kopplas bort från den regionala livsuppehållande apparaten .
Det är viktigt att fastställa de kunskaper och möjligheter som finns i våra regioner inom den högteknologiska sektorn .
Det är särskilt viktigt mot bakgrund av rapporterna i media som säger att Europa snabbt håller på att tappa mark till Förenta staterna i de framtida högteknologiska tillväxtbranscherna .
Verksamheten inom den förra programrundan visar också på ett tydligt sätt vad riktlinjer inte skall handla om .
De skall inte handla om att skapa ytterligare byråkrati och snåriga bestämmelser .
De skall inte handla om att ändra inriktning och politik när man kommit halvvägs genom projektet , vilket resulterar i oundvikliga förseningar och outnyttjade medel , i synnerhet mot bakgrund av det nya budgetkravet .
Tillämpningen och genomförandet av riktlinjerna kan inte överlåtas till personlig tolkning av någon tjänsteman vid kommissionen eller den nationella statliga förvaltningen .
Det måste råda en intern sammanhållning vid kommissionsdirektoratet , samtidigt som man respekterar de specifika lokala och regionala aspekterna av kommissionens program .
Slutsatsen blir att vi måste se till att riktlinjerna blir breda , vägledande och flexibla för att hjälpa våra programansvariga och de som tar emot medel , och att erhålla maximala möjligheter från våra nya förnyelseområden .
Om vi kan tillföra en anda av entreprenörskap i våra fattiga och strukturellt svaga regioner , kommer vi till sist att få dem på rätt köl när det gäller att dra till sig större volymer investeringskapital , som kommer att vara nyckeln till framgång .
Det är så vi skall bedöma hur framgångsrika dessa riktlinjer blir : Om EU : s regionalpolitik med bra , gedigna och kreativa riktlinjer kan skapa nya möjligheter och göra det möjligt för våra fattiga och strukturellt svaga regioner att efter förmåga bidra till EU : s framtida tillväxt och välstånd .
Herr talman , herr kommissionär , bästa kolleger !
Jag vill tacka Schroedter för ett bra betänkande .
Hon har med omsorg satt sig in i ärendet och under utskottsbehandlingen på ett bra sätt beaktat de många ändringar som gjorts i detta betänkande .
Föredraganden har också helt riktigt konstaterat att parlamentet inte i tid hörts angående riktlinjerna .
Nu är man mycket försenad i frågan .
Förhoppningsvis hjälper dock parlamentets ställningstaganden till vid bedömningen av programmen efter halva vägen och vid det praktiska genomförandet av dem .
Med tanke på tidpunkten har betänkandet under behandlingen blivit alltför omfattande .
Man har där samlat detaljerade frågor och till och med sådant som redan tagits upp i tidigare betänkanden .
I detta skede är det viktigare att koncentrera sig på att bedöma på vilket sätt man genom den här processen skulle kunna styra unionens regionalpolitik med tanke på att målet är att minska den regionala obalansen .
Vår grupp framhåller subsidiaritetsprincipen , medlemsstaternas ansvar och de lokala aktörernas roll vid utarbetandet och genomförandet av programmen .
Det är speciellt viktigt att involvera de små och medelstora företagen i planeringen och genomförandet av programmen .
Vår grupp anser det också vara viktigt att ta mer hänsyn till utomeuropeiska områden och andra ytterområden och vi vill öka växelverkan mellan städerna och landsbygden .
Vi motsätter oss ett alltför långtgående förmyndarskap från unionens och medlemsstaternas centralförvaltningars sida och kräver att den byråkrati som fått fotfäste vid utarbetandet och genomförandet av programmen bantas ned .
Effekten av projekt som genomförts med hjälp av unionens bidrag har alltför ofta försvagats på grund av långsamt beslutsfattande och krånglig förvaltning .
Ofta har man beviljat anslag till projekt som inte gett regionen någon bestående nytta .
Projekten måste bli effektivare , mer flexibla och de måste leda till bättre resultat .
I samband med utarbetandet av betänkandet fördes det också en intressant debatt om unionens regionalpolitik i största allmänhet .
Det var första gången för oss nya ledamöter och detta är en mycket intressant process .
Detta är ett bra betänkande , vår grupp ställer sig bakom det .
Herr talman , herr kommissionär , ärade ledamöter !
Som ett bevis på att detta parlament ännu inte har kommit över sin roll som rådgivande och underordnad institution , är det utmärkta betänkandet från min gruppkollega Elisabeth Schroedter ännu inte framlagt i kammaren på grund av att planerna för den regionala utvecklingen under tiden 2000-2006 för mål 1-områden redan har legat flera månader på kommissionens sekretariat .
Med hänsyn till detta måste detta parlament hur som helst , innan det godkänner gemenskapens stödramar för den period det gäller , kräva att dessa analyseras och debatteras i kammaren i ljuset av just de inriktningar vi lägger fram i dag , där vi särskilt trycker på deras förmåga att skapa sysselsättning i de fattigaste eller minst utvecklade områdena , och att vi därigenom bidrar till att förändra de nuvarande negativa tendenserna till ojämlikhet i det europeiska samhället och arbetar för ett rättvisare Europa .
Herr talman !
Vi får inte glömma bort att det främsta strategiska målet med strukturfonderna och Sammanhållningsfonden och samordningen av dessa är att uppnå en ekonomisk och social sammanhållning .
Vi är skyldiga att medverka till utformandet av riktlinjerna och även i utvärderingen av resultaten .
Och detta för att vi är medborgarnas företrädare i medborgarnas Europa , och inte bara i ett staternas och regionernas Europa .
Vi kan konstatera att fonderna är en nödvändig , men otillräcklig förutsättning för att uppnå ekonomisk och social sammanhållning .
Om vi använder oss av bruttonationalprodukten per invånare som den enda indikatorn kan vi missta oss .
Några av kollegerna har redan talat om arbetslösheten , om nedgången i demografin .
Vi borde undersöka ett antal indikatorer som tillåter oss att bedöma situationen och utvecklingen i sådana regionala samhällen där situationen är värre än i de övriga .
Av vissa av de betänkanden som i dag har lagts fram inför parlamentets plenum framgår det att arbetslösheten i de 25 mest framgångsrika europeiska regionerna är fem gånger lägre än i de 25 minst framgångsrika regionerna .
Det tvingar Europaparlamentet , herr kommissionären och kommissionen att agera på ett beslutsamt och strategiskt sätt .
Jag håller med om att Europaparlamentet inte hade någon möjlighet - eller inte fick någon sådan för att mandatperioden snart skulle vara över - att diskutera dessa riktlinjer .
Men jag tror inte att betänkandet kommer att dröja .
Vi behöver tillsammans fundera över hur de nya programmen med mål 1 och de planer för regional utveckling som har utvecklats innan riktlinjerna träder i kraft , skall kunna bli föremål för en granskning och en riktig utvärdering .
Det krävs en samordning av programmen med de olika målen .
Vi ställer alla kravet att även parlamentet , när halva verksamhetstiden för programmen har gått och det är dags att utvärdera riktlinjerna , skall inta en ledande roll , för vi är medborgarnas företrädare .
Medborgarna kan inte acceptera att Europeiska unionen fattar beslut på ett så till synes byråkratiskt sätt .
De förväntar sig att den politiska dimensionen finns med , att man visar ansvar , att det finns en kommunikation med medborgarna .
Det är det vi i dag vill be herr kommissionären om .
Jag hoppas att han , efter sina senaste erfarenheter som regional ordförande , kommer att gå med på att föreslå vissa indikatorer och en strategi till förmån för den ekonomiska och sociala sammanhållningen och inte bara för produktiviteten .
Herr talman !
Jag stöder huvudförslagen i betänkandet rörande förvaltningen av strukturfonderna och Sammanhållningsfonden för perioden 2000-2006 och betänkandets huvudrekommendationer vilka inkluderar följande : Det måste alltid råda ett samordnat förhållningssätt till finansieringen ur EU : s strukturfonder och Sammanhållningsfonden .
Detta innebär att det måste råda ett heltäckande partnerskap mellan lokala myndigheter och nationella regeringar med hänsyn till hur dessa medel skall användas .
Medlemsstaterna uppmanas att lägga större vikt vid samordnade strategier för en förnyelse av förhållandena mellan städer och landsbygd .
Denna senare fråga är av särskild betydelse .
Samtidigt som förnyelsen av våra stadsområden är mycket viktig måste vi alltid hitta en balans i vår politik mellan främjandet av landsbygdens utveckling och förbättringen av livskvaliteten för dem som bor i städerna .
Vi har inte för avsikt att bygga ett Europa som bara består av städer .
Strukturfonderna har spelat en viktig roll för utvecklingen av både städer och landsbygd i perifera länder , huvudsakligen genom förbättring av vägar , vattenrening och transportnät som har samband med detta .
Denna process kommer att fortsätta i överensstämmelse med riktlinjerna för finansiella utgifter , vilka fastställdes av EU : s politiska ledare vid toppmötet i Berlin förra året , och vilka stöddes av parlamentet vid dess sammanträdesperiod i maj .
Tongivande EU-program mellan 1989 , 1993 , 1994 och 1999 har verkligen hjälpt till att förbättra den ekonomiska konkurrenskraften i perifera länder och mål 1-regioner i Europeiska unionen .
Det viktiga är nu att konsolidera och befästa de framsteg som gjorts hittills .
Detta kommer att garantera att randområdena och de yttersta randområdena , de fattigare regionerna i Europeiska unionen , hamnar i en ställning där de kan nå framgångar inom det nya euroområdet , såväl som inom den ständigt expanderande inre marknaden där det råder fri rörlighet för varor , personer , tjänster och kapital .
Sammanfattningsvis - medan viktiga infrastrukturprojekt fått medel från Europeiska regionala utvecklingsfonden och Sammanhållningsfonden , bör vi komma ihåg att Europeiska socialfonden har spelat en mycket viktig roll vad gäller hjälp till de fattiga i samhället .
Socialfonden har verkligen förbättrat våra institutioner för högre utbildning , finansierat våra studieprogram för personer som redan innehar examensbevis och fått till stånd omfattande program som syftar till att bekämpa ungdoms- och långtidsarbetslöshet , hjälpa personer som lämnat skolan vid ett tidigt skede och främja en högre standard vad gäller läskunnigheten hos vuxna .
Herr talman !
Jag har tidigare flera gånger varit oense med föredraganden , när det gäller regionalpolitiska frågor , men denna gång delar jag hennes uppfattning .
Jag vet inte om detta uppmuntrar henne att fortsätta i samma riktning , men i vilket fall som helst skulle jag vilja framföra mina gratulationer .
Den andra punkten som jag skulle vilja ta upp är det önskemål som McCarthy och jag framförde i egenskap av föredraganden för den allmänna förordningen .
Jag skulle alltså föredra att riktlinjerna fogades till förordningen som bilaga .
Detta har tyvärr inte skett , och den som bär ansvaret för detta är inte Bernié utan det förutvarande utskottet .
Jag framför detta för att upprepa parlamentets ståndpunkt .
Den tredje punkten som jag skulle vilja ta upp är att jag stöder riktlinjerna i stora drag , i den mån de inte avviker från de anmärkningar vi gjort .
Riktlinjerna är till stor hjälp för medlemsstaterna , jag vill särskilt framhålla hur stor betydelse kommissionen tillmäter frågan om hållbar utveckling och ökad sysselsättning , i synnerhet när det gäller likvärdiga möjligheter och transportfrågor .
Detta kan åtminstone jag personligen helt och hållet instämma i .
Sedan skulle jag i egenskap av öbo vilja kritisera att man försummat frågan om öarnas utveckling .
Man lägger inte tillräckligt stor vikt vid detta , och det är heller inte första gången .
Under mina fem år som ledamot av parlamentet har jag upprepade gånger berört denna fråga .
Herr kommissionär , jag kommer även i fortsättningen att ta upp denna fråga , för i artikel 158.1 i Amsterdamfördraget finns en bestämmelse som handlar om en helhetspolitik för öarna .
Följaktligen borde kommissionen nu äntligen ta och granska den konkreta frågan .
Sedan , herr kommissionär , är det nu äntligen dags att genomföra programmen , även medlemsstaterna måste alltså ta sitt ansvar och sköta sina uppgifter på ett riktigt sätt .
Beträffande oss här i parlamentet vill jag påminna om att det finns en uppförandekod för relationerna mellan parlamentet och kommissionen , som undertecknades i maj .
Jag är förvissad om att denna kod kommer att följas och att parlamentet kommer att hållas underrättat om detaljer i fråga om genomförandet av programmen .
Herr talman , herr kommissionär , kära kolleger !
Under den en och en halv minut jag har till mitt förfogande skulle jag till att börja med vilja lyckönska kollegan Schroedter .
Jag tror att många redan gjort det , men jag tycker att hon förtjänar det eftersom hon varit mycket öppen och lyhörd för förslag från andra och jag tror att det är tack vare hennes tillgänglighet som betänkandet blivit så bra .
Jag instämmer i hennes beklagande över att parlamentet på sätt och vis hoppat på tåget i farten när det gäller riktlinjerna , eftersom förhandlingsförfarandet med staterna i dag har kommit så långt att det är svårt att tro att detta betänkande får någon direkt inverkan , vilket jag beklagar .
Det förefaller därför som om man i betänkandet behöver föregripa och fastställa riktlinjerna för revideringen efter halva tiden år 2003 , och även påverka den andra delen av programmen efter 2003 .
Jag skulle kort sagt vilja säga att vi går in i en förvaltningsperiod för programplaneringen 2000-2006 , som inte får vara en rutinperiod , av den enkla anledningen att vi står inför två stora utmaningar .
Den första gäller harmoniseringen av politiken för den nationella fysiska planeringen och politiken för regional utveckling .
Anslagen räcker inte till för att bedriva utveckling , när det finns brister i infrastruktur eller offentlig service .
Det är alltså en grundläggande fråga vi måste ställa oss : hur kan vi se till att unionens politik flätas samman med den extra nationella politiken för fysisk planering .
Den andra utmaningen handlar om utvidgningen , som naturligtvis får avsevärda konsekvenser såväl på budgetområdet som geografiskt .
Detta är två uppgifter som jag uppmanar kommissionären att genomföra och där jag ber honom att ta med oss i diskussionerna .
I denna tid av naturkatastrofer skulle jag ändå vilja ta upp frågan om strukturfondernas utnyttjande .
Vi vet att det åligger varje stat att fördela en del av totalanslaget .
Det får inte bli så som staterna har en tendens att vilja , att Europa försvinner helt .
I dag anklagar den allmänna opinionen och pressen oss för att vara otillgängliga medan vi skall finansiera en stor del av de nationella ansträngningarna .
Jag tror att vi måste kunna säga det högt och tydligt .
Jag tror att vi också måste inrätta eller be medlemsstaterna att ansvara för information om det europeiska stödet varje gång det utnyttjas för att reparera skador som orsakats av naturkatastrofer eller olyckor .
Herr talman !
Prioriteringen av ekonomiska kriterier och monetära kriterier ökar orättvisorna i alla dess former .
För den franska planens experter exempelvis är det mest troliga scenariot i dag att de regionala skillnaderna ökar i varje land .
Men strukturfonderna har bidragit till att bromsa denna process .
Vårt projekt med ett Europa som kan uppfylla sociala behov syftar till att höja levnadsstandarden och göra den enhetlig .
Genomförandet skulle sannolikt leda till att sådana fördelningsinstrument som strukturfonderna skulle utvidgas .
Vi föreslår framför allt en enhetlig kapitalskatt , som skulle göra det möjligt att bidra till fonder som kan åtfölja harmoniseringen av socialförsäkringssystemen och en minskning av arbetstiden på europeisk nivå .
Men när kommissionen ombeds att lägga fram riktlinjer gör den det med ett beklagande och på ett luddigt sätt .
Det betänkande som i dag läggs fram ger på nytt politiken en plats .
Det är ett steg på väg mot en hållbar politik för sysselsättning och utveckling .
Och det är det som gör att vi kan rösta för den .
Herr talman !
Även jag vill tacka föredraganden för ett utmärkt arbete .
Mer än någonsin tidigare kommer Europa under de kommande åren , på grund av den utmaning som globaliseringen och östutvidgningen medför , att behöva klara och tydliga riktlinjer när det gäller program för att åter få fart på den ekonomiska utvecklingen .
I det avseendet måste Europa som helhet , och varje enskild medlemsstat , på bästa sätt utnyttja alla sina resurser och möjligheter , och därmed också de strukturfonder som är tillgängliga .
För att göra det krävs en europeisk kommission som , utöver de goda avsikterna , är tydligare i sina riktlinjer och anstränger sig maximalt i arbetet att kontrollera hur medlemsstaterna utnyttjar dessa resurser .
Italien till exempel har under de senaste åren haft problem när det gällt att utnyttja strukturfonderna , framför allt på grund av en överdriven byråkrati , bristfällig information och ett bristande engagemang från de ekonomiska och sociala operatörerna på lokal nivå .
Det är därför i första hand två punkter jag vill rikta kommissionens uppmärksamhet på : för det första gäller det att på bästa sätt utnyttja samråd som en metod att samordna lokala och regionala operatörer och göra dem delaktiga i besluten , just för att undvika obalanser och orättvisor .
För det andra måste de administrativa processerna förenklas och göras mer lättillgängliga , eftersom de alltför ofta blir onödigt långa och komplexa , till den grad att de äventyrar tillgången till fonderna , något som framför allt de små och medelstora europeiska företagen klagar över .
Herr talman !
Låt mig avslutningsvis säga att det är ganska allvarligt att kommissionen i sitt meddelande bara ägnar bristfällig uppmärksamhet åt de territoriella avtalen och framför allt kampen mot arbetslösheten vad gäller kvinnor och ungdomar .
Herr talman !
I likhet med min kollega Evans , tycker jag att det är synnerligen trevligt att stiga upp i talarstolen och hålla mitt första tal i denna kammare om denna mycket viktiga fråga , särskilt på grund av att jag företräder en del av Förenade kungariket , West Midlands , som hittills dragit nytta av i synnerhet finansiering från mål 2 .
Men det betänkande som behandlas i kammaren i kväll är ett utmärkt exempel på - om vi inte är väldigt försiktiga - hur vi kan lägga fram mycket storslagna idéer som saknar det innehåll som gör dem relevanta för de personer som direkt drar nytta av dem .
Betänkandet i sig självt har ett gott syfte men , som så ofta när vi behandlar dessa frågor , saknar ett tydligt syfte och en sund verksamhetsbas .
Detta är skälet till varför jag och min grupp lägger fram tre viktiga ändringsförslag och tillägg till texten - inte för att ta bort något från förslaget , utan för att göra det mer relevant för de som det är avsett att ge vägledning .
Låt mig förklara hur vi har tänkt här .
För det första vill vi se till att strukturfonderna och Sammanhållningsfonden används på ett lämpligt sätt .
Erfarenheten visar , i egenskap av företrädare för skattebetalarna i Europeiska unionen , att vi bör - att vi måste - kräva finansiell redlighet och öppenhet i samband med utbetalningarna och kontrollen av dessa pengar .
Våra ändringsförslag och tillägg har därför att göra med uppfyllandet av vad som är känt som " valuta för pengarna " indikatorer under förfarandet där beviljande av anslag sker .
Vi får dessutom alltför ofta se att enorma belopp används inom projekt vars resultat man vet kommer att bli otydliga redan vid början av programperioden .
Men halvvägs igenom eller vid slutet av denna period finns det inget effektivt sätt att avsluta projektet på , om det inte visat sig vara framgångsrikt .
I våra tillägg uppmanar vi därför till att man skall skapa bestämmelser om strategier för ett praktiskt genomförbart avslutande , så att vi inte bara kan få den nödvändiga garantin mot fortgående kostnader som ofta skattebetalarna får står för , utan så att vi också kan undvika det väl inövade syndromet som innebär att vi offrar ytterligare pengar på ett hopplöst projekt .
Slutligen efterlyser vi en förändring vad gäller den balans och den metod som används vid utbetalningen av medel .
Det bör vara ett större deltagande från den privata sektorns sida , vilket kommer att ge realistiska ekonomiska perspektiv vid utarbetandet av finansieringsplanerna .
Dessutom måste de finansierade projekten - i stället för att vara småskaliga , intäktsbaserade projekt , vilka är svåra att övervaka - bli mer storskaliga , eftersom de positiva effekterna då blir mer uppenbara .
På så sätt kommer det ofta utbasunerade behovet av öppenhet i samband med användningen av dessa medel att minska , och det kommer också frestelsen att i det längre perspektivet på ett onödigt sätt förlita sig på den lokala skattebasen i områden där projekten genomförs .
Europaparlamentet kommer sålunda att visa hur allvarligt man ser på behovet av sådana reformer .
Om dessa ändringar av betänkandet stöds av kammaren i dag , menar jag att detta kommer att förflytta oss till nästa fas , då vi kan åstadkomma de historiska mål som fonderna syftar till , dvs. att på ett ekonomiskt hållbart sätt hjälpa medborgarna i de eftersatta områdena i Europeiska unionen att få en tillfredsställande levnadsstandard ; inte genom att ge allmosor , utan att ge hjälp till självhjälp .
Jag uppmanar kammaren att stödja dessa ändringsförslag .
Herr talman , herr kommissionär , värderade kolleger !
Även jag skulle vilja gratulera föredraganden och tacka henne för hennes stora och seriösa arbetsinsats .
Det råder inget tvivel om att Europeiska unionens strukturpolitik och sammanhållningspolitik är de viktigaste instrumenten för att skapa förutsättningar för utveckling och för att minska de ekonomiska och sociala klyftorna mellan regionerna .
Trots de åtgärder som vidtagits består dessa klyftor , och i synnerhet när det gäller arbetslösheten är de mycket större än man kan acceptera .
För att denna politiks mål skall uppnås i största möjliga utsträckning är det nödvändigt att de politiska insatserna samordnas och att de organiseras med ledning av väl genomtänkta , jag skulle vilja säga intelligenta , riktlinjer .
Vi får inte glömma att dessa politiska insatser , när de är effektiva , är synliga också för de europeiska medborgarna , som drar nytta av dem och som ser en direkt förbättring av sin livskvalitet .
Vi får inte glömma att man särskilt måste uppmärksamma Europeiska unionens avsides belägna regioner och dess öregioner , för deras geografiska läge medför stora hinder för deras ekonomiska och sociala utveckling , såvida inte kommissionen kanske har för avsikt att bygga broar eller tunnlar för att förbinda öarna med det europeiska fastlandet .
Avslutningsvis skulle jag vilja framhålla att strukturpolitiken i sin helhet måste bli mera flexibel , så att den anpassas till föränderliga situationer och därigenom bättre kan möta de nya utmaningar och nya möjligheter , som uppstår när vi nu har gått in i ett nytt millennium som vi alla knyter varma förhoppningar till .
Herr talman !
Schroedters betänkande innehåller utan tvivel ganska många viktiga iakttagelser , och därför vill jag gratulera henne .
Jag anser emellertid att vi borde hysa ännu större oro när det gäller gemenskapens regionalpolitik , dess inriktning och effektivitet .
Man kan sammanfattningsvis konstatera att den enorma massarbetslösheten långt ifrån att lindras tvärtom förvärras ytterligare genom strukturpolitiken .
Jordbruksekonomin och jordbruksregionerna drabbas ohjälpligt av den regionalpolitik som bedrivs , med dramatiska följder för sysselsättningen på landsbygden och för jordbrukarnas levnadsvillkor , framför allt i södra Europa .
Den regionala obalansen ökar dramatiskt inom medlemsstaterna .
Om vi betraktar uppgifterna i den sjätte rapporten , skall vi finna att den regionala obalansen har ökat enormt under de senaste tio åren .
Man uppmärksammar nästan inte alls de enorma problemen i unionens öregioner , där bristerna i fråga om infrastruktur , transporter , kommunikationer och energi leder till en ständigt fortgående avfolkning .
Ansvaret för detta bärs såväl av unionens regionalpolitik som av dess ekonomiska och sociala politik över huvud taget .
Stora delar av Europas befolkning fördömer skarpt denna politik som farlig och antifolklig .
De nya riktlinjerna har tyvärr samma inriktning , och det finns ingenting som tyder på att inriktningen kan förändras genom att man tillämpar dessa riktlinjer .
Herr talman , kära kolleger !
Låt mig säga några korta ord för att betona två punkter , som dessa betänkanden påminner oss om , och som har en strategisk betydelse för det perspektiv vi har på unionen .
Den första är den väsentliga och centrala betydelse som vi fortfarande fäster vid den ekonomiska och sociala sammanhållningen .
Vi oroar oss också över nyheter om att kommissionens känsla för betydelsen av detta mål avtar .
Vi kommer att fortsätta att betrakta unionens ekonomiska och sociala sammanhållning som central .
För det andra håller jag med om de ord vi här har hört från en kollega angående öarna , och jag vill även uppmärksamma regionerna i gemenskapens yttersta randområden .
Vi skulle i framtiden vilja se mer djärvhet i hanteringen av regionerna i de yttersta randområdena , som beträffande mitt land när det gäller Azorerna och Madeira .
Jag vill passa på detta tillfälle att fråga om kommissionen skulle kunna redogöra för skälen till att kommissionens rapport om gemenskapens yttersta randområden , som parlamentet har väntat länge på , är försenad ?
Herr talman !
Först vill jag tacka föredraganden , också för hennes beredvillighet att ta med synpunkterna från vår sida i betänkandet .
Herr talman , mina damer och herrar , herr kommissionär !
Med hjälp av riktlinjer skall medlemsstaterna erbjudas en orientering i att uppnå reformmålen inom ramen för programmeringen .
Här resulterar dock kommissionens direktiv , tvärtemot anspråken på att vilja erbjuda en orientering , snarare i en anbudskatalog över möjliga åtgärder inom de olika politiska fälten .
Ändå är den egentliga avsikten att ange riktning och visa på vad som bör prioriteras .
Jag delar helt föredragandens åsikt om att kommissionens dokument tyvärr innehåller för få rekommendationer till medlemsstaterna när det gäller förenkling av förvaltningsförfarandet , och jag vill understryka krav som att förhandlingarna koncentreras till att främja en gynnsam miljö för arbetsintensiva små och medelstora företag , en tydlig målsättning för alternativa finansieringskällor inklusive bestämmelser för riskkapital och privat finansiering , starthjälp för företag inklusive ny informationsteknik liksom investeringar på innovativa områden .
Särskilt stöd vill jag ge åt ett ändringsförslag från min grupp under siffran 10 , vilket skall garantera att den privata sektorn i rimlig utsträckning inkluderas i planeringen och genomförandet av projekten .
Fru Schroedter , jag skulle uppskatta om ni , inte minst med tanke på subsidiaritetsprincipen , ville ta med detta ändringsförslag i era positiva överväganden .
Herr talman , herr kommissionär !
I utskottet för sysselsättning och socialfrågor var vi eniga om kravet på att det viktigaste och strategiskt korrekta var att stödja strukturfondernas och Sammanhållningsfondens insatser för en ökad sysselsättning bland de arbetslösa och för jämlikhet mellan kvinnor och män .
Tyvärr har inte det kravet beaktats i Schroedters utmärkta betänkande , trots att det finns många bevis - något som vi senare kommer att få se i Berends betänkande - på hur dessa fonder på ett fantastiskt sätt stöder de sämst utvecklade regionerna att överbrygga det avstånd som skiljer dem från de mest välutvecklade regionerna i Europa .
Dessa regioner håller på att expandera , vad BNI beträffar .
De håller på att expandera i konkurrenskraft , men inte alla får ta del av den ökade rikedomen , för det är inte sysselsättningen som ökar , och skillnaderna i de olika regionerna beträffande arbetstillfällena kvarstår .
Herr kommissionär , läs yttrandet från utskottet för sysselsättning och socialfrågor och prioritera detta , för det är där det stora problemet för medborgarna ligger .
Och var strategisk i samband med granskningen och beviljandet av fondmedel , och ta hänsyn till behovet av sysselsättning , för det är definitivt något som strukturfonderna och Sammanhållningsfonden kräver .
Herr talman !
Riktlinjerna måste på ett korrekt sätt kunna styra och effektivisera programmen under den avgörande sjuårsperioden 2000-2006 , så att man äntligen kan förverkliga hållbar utveckling och förbättrad sysselsättning , i synnerhet bland kvinnor och ungdomar , och så att man kan åstadkomma balans mellan miljöpolitiken och den ekonomiska och sociala politiken .
Det är särskilt viktigt att ta itu med städernas växande problem , att bibehålla arbetstillfällena på landsbygden , att stödja jordbruksregionerna och , naturligtvis , att erbjuda likvärdiga utvecklingsmöjligheter för Europeiska unionens öar och för de grekiska öarna , som utgör hälften av unionens öar , allt i enlighet med artikel 158 i fördraget .
Sammanhållningspolitiken måste stärkas ytterligare , för ett Europa med enorma klyftor i fråga om levnadsstandard i olika regioner kan inte vara vare sig trovärdigt eller livskraftigt . .
( FR ) Herr talman , mina damer och herrar parlamentsledamöter !
Det var mycket intressant att noga lyssna till kommentarerna , som ibland var kritiska , och förslagen nyss i era inlägg med utgångspunkt från Schroedters betänkande .
Fru föredragande , mina damer och herrar !
Alla förstår anledningarna , tidsfristerna - jag skall snart återkomma dit , - och vilka dessa tidsfrister och förseningar än må vara , eftersom det är nu som vi diskuterar detta betänkande , anser jag för kommissionens räkning , att det kommer vid rätt tillfälle , det gäller ju riktlinjerna för 2000-2006 , för det är ju nu som vi skall inleda den nya programplaneringsperioden för regionalpolitiken .
Fru föredragande !
Ni erinrade med rätta om att även om det faktiskt huvudsakligen åligger medlemsstaterna och regionerna att fastställa sina egna prioriteringar när det gäller utveckling , kräver och motiverar Europeiska unionens medfinansiering av programmen att man också beaktar gemenskapens prioriteringar , så som de diskuterats och godkänts här , för att främja denna gemenskapsdimension av den ekonomiska och sociala sammanhållningen , som många av er erinrat om med kraft .
Mina damer och herrar !
Jag skulle också ha önskat att om en stund återkomma till riktlinjernas roll och struktur innan jag tar upp de huvudsakliga kommentarerna eller kritiska åsikterna som ni , fru föredragande , eller ni själva , mina damer och herrar , har framfört .
När det gäller riktlinjernas roll och struktur erinrade ordförande Hatzidakis , föredraganden och McCarthy om att dessa riktlinjer har till uppgift att hjälpa de nationella och regionala myndigheterna med att förbereda sin programplaneringsstrategi för vart och ett av målen 1 , 2 och 3 inom strukturfonderna , liksom deras förbindelser med Sammanhållningsfonden .
Det handlar om att lägga fram kommissionens prioriteringar med stöd av tidigare erfarenheter från att genomföra programmen , likaväl som nuvarande gemenskapspolitik knuten till ingripanden genom strukturfonderna .
Och målsättningen är just att dessa prioriteringar skall bidra till ett bättre utnyttjande , ett optimalt och effektivt utnyttjande av gemenskapsåtgärderna , inbegripet , herr Bradbourn , att vid rätt tillfälle utnyttja prestandareserven vars mål bl.a. är att uppmuntra till ett optimalt och effektivt utnyttjande av de offentliga europeiska medlen .
Och när jag talar om optimalt utnyttjande menar jag såväl på nationell nivå som regional nivå .
Herr Seppänen !
Jag nämner därför också - när vi talar om den nationella nivån - kopplingen till Sammanhållningsfonden .
Så långt målsättningen med dessa riktlinjer .
När det gäller innehållet rör det sig som ni vet , mina damer och herrar parlamentsledamöter , om tre strategiska prioriteringar som er föredragande mycket tydligt och samtidigt mycket ivrigt , förstod jag av anförandet nyss , erinrat om .
Den första prioriteringen gäller förbättrad konkurrenskraft för de regionala ekonomierna för att inom alla sektorer , men särskilt inom den privata sektorn , såsom Berend sade , skapa så många seriösa , starka och beständiga arbetstillfällen som möjligt .
Konkurrenskraft för de regionala ekonomierna , för alla regionala ekonomier och särskilt , herr Evans , för Wales , men inte bara Wales .
Och eftersom flera av er på nytt betonat något som föreföll vara bortglömt skall jag tillägga de regionala ekonomierna i de europeiska regioner som hindras av det faktum att de ligger långt bort , vare sig det gäller perifera områden , öregionerna eller , naturligtvis , de yttersta randområdena som ligger allra längst bort .
Kanske kan jag i det sammanhanget säga till Ribeiro i Castro som ställt frågan till mig att , såsom jag skrivit till presidenterna i vart och ett av dessa yttersta randområden , har kommissionen begärt ytterligare litet tid för att offentliggöra den rapport som förväntas av den .
Vi fick när det gäller de yttersta randområdena skrivelserna från de olika regeringarna ganska sent , men det behöver inte vara en ursäkt , bara en förklaring .
Vi måste alltså beakta dessa skrivelser och utföra detta mycket viktiga arbete .
Jag deltog personligen i ett möte med företrädare för de yttersta randområdena den 23 november och vi ansåg inom kollegiet att vi behövde ytterligare några veckor för att åstadkomma en rapport som är i nivå med de mycket seriösa och allvarliga problemen och förväntningarna från dessa yttersta randområden , och jag tackar för att ni har förståelse för detta .
Så långt den första prioriteringen , nämligen de regionala ekonomiernas konkurrenskraft .
Den andra prioriteringen som flera av er betonat - särskilt Puerta , men även andra - jag gör ingen inbördes prioritering dem emellan , handlar om att stärka den sociala sammanhållningen och sysselsättningen , särskilt genom att på ett bättre sätt än tidigare uppvärdera de mänskliga resurserna .
Mina damer och herrar parlamentsledamöter !
En europeisk union med färre skillnader mellan länderna , vilket för övrigt bevisar att Sammanhållningsfonden är effektiv och gör nytta , men där man samtidigt när det gäller arbetslösheten konstaterar - ni skrev det fru talman - att skillnaderna ökar mellan de 15 eller 20 rikaste regionerna och de 15 eller 20 fattigaste , eller de sämst lottade , är en situation som är , som skulle vara , omotiverad och oacceptabel .
När det gäller mig själv - med tanke framför allt på att jag håller på att sätta mig in i den europeiska integrationen och den regionala utvecklingspolitiken , - är det en situation som jag inte kan acceptera och jag har för avsikt att så långt det är möjligt och med ert stöd ställa anslag som jag ansvarar för till förfogande för denna förbättrade sociala , mänskliga , territoriella sammanhållning , bl.a. för att vi inte skall få ett Europa med två hastigheter , ett Europa med flotta kvarter och ett annat med fattiga förorter , något som jag tidigare talat om .
Den tredje målsättningen gäller utvecklingen i städerna och på landsbygden , inom ramen för en rättvis territorialpolitik .
I riktlinjerna tas hänsyn till två horisontella principer : landsbygdsutveckling och , fru föredragande , jag innefattar i landsbygdsutveckling också frågan om hållbara transporter som jag personligen fäster stor betydelse vid sedan länge - bl.a. när jag tänker på min tid som miljöminister i mitt land - och den andra principen handlar om lika möjligheter , framför allt för män och kvinnor , liksom den europeiska strategin för sysselsättning och ramen för den ekonomiska och monetära unionen .
Avslutningsvis och för att bemöta den oro ni uttryckt - och särskilt ni , fru föredragande - erinras i dessa riktlinjer om betydelsen och definitionen av integrerade strategier för utveckling eller omställning , som bland alla dessa prioriteringar ger den största chansen till synergier , till åtgärder och till att inrätta ett decentraliserat partnerskap .
Ni oroade er för vad som skulle kunna framstå som avsaknad av hänvisning till detta partnerskap - det nämns ändå tydligt på sidan 5 i dessa riktlinjer , men jag vill gärna erinra om det - eftersom ni ber om det - att för mig är detta partnerskap - och jag har varit ansvarig tillräckligt länge för en region i mitt land för att kunna säga det ärligt - ett verktyg , det är hävstångseffekten av lokal intelligens , vare sig den finns inom den offentliga sektorn , de folkvalda , den sociala sektorn och undervisningssektorn , föreningarna eller den privata sektorn .
Ett decentraliserat partnerskap , och jag vill i detta sammanhang för att svara Angelilli naturligtvis ta upp de territoriella pakterna , som är en av möjligheterna inom detta decentraliserade partnerskap .
Detta var anledningarna till att riktlinjerna presenterats efter prioriteringar per område , eftersom de måste beaktas på olika nivåer utifrån varje medlemsstat och regions särskilda situation , i enlighet med respektive målsättning .
Jag skulle nu snabbt vilja kommentera några av era anmärkningar , mina damer och herrar , till att börja med om förfarandet .
Det stämmer att kammaren tillfrågades sent .
Tillåt mig erinra om att när riktlinjerna antogs av kommissionen , i form av ett förslag i februari 1999 , efter ett nytt förfarande som skulle underlätta framläggandet av kommentarer om texten , överlämnades de omedelbart till parlamentet av min företrädare , Monica Wulf-Mathies .
Men med tanke på det nära förestående valet till Europaparlamentet var det först efter att texten definitivt antagits , i juli 1999 , som kammaren kunde börja granska dessa riktlinjer .
När jag nu befinner mig bland er , mina damer och herrar , vill jag försäkra er om att i förhandlingarna om programmen , som precis bara har börjat för de flesta medlemsstater - ordförande Hatzidakis frågade mig om det - kommer era kommentarer absolut att beaktas .
Och jag kan dessutom försäkra er om att när kommissionen antar riktlinjerna inför det som kallas översyn efter halva tiden , såsom arbetsordningen föreskriver , kommer man också att beakta kammarens uppfattning , vilken uttrycks i betänkandet .
När det sedan gäller sakfrågan , riktlinjernas roll , fru föredragande , betonade ni att det är just inom denna ram som det gäller att tillhandahålla riktlinjer om ett antal europeiska målsättningar , som ofta är mycket precisa .
Jag skall bara nämna några : genomförande av en politik inom olika sektorer , bättre utnyttjande av offentliga medel , stöd till de olika parterna för att gemensamt utarbeta regionala eller nationella programplaneringar , etc .
Kommissionen noterar detta , men flera av dessa riktlinjer eller dessa frågor faller snarare under andra dokument , såsom Vademecum eller dokumentet om arbetsmetoder .
Jag skulle avslutningsvis vilja inrikta mig på vissa frågor ni tagit upp , fru föredragande .
Jag tänker exempelvis på idén att riktlinjerna inte är tillräckligt specifika när det gäller rekommendationerna .
Detta påstående i ert betänkande måste ses i sammanhanget med förhandlingarna förra våren .
Kommissionen höll sig till texten i artikel 10 i den allmänna förordningen om strukturfonderna , där det anges att dessa riktlinjer skall ge medlemsstaterna allmänna vägledande riktlinjer , som bygger på relevant och överenskommen gemenskapspolitik .
Det är själva texten jag citerat , inom citationstecken .
Riktlinjerna kan inte ersätta programplaneringen eller ex ante-utvärderingarna som måste vara det instrument som kan ange prioriteringarna och effektiviteten i dessa program .
Fru föredragande !
Ni tog sedan upp avsnittet med riktlinjer för utveckling av stadsmiljön och landsbygden och ansåg att utvecklingen av stadsmiljön inte beaktats tillräckligt .
Tvärtom , tycker jag .
Jag vill framhålla att kommissionen fäster stor betydelse , även i framtiden , vid stadsmiljön inom sammanhållningspolitiken .
Jag hade för övrigt tillfälle att säga det till samtliga ministrar med ansvar för stadspolitiken vid ett möte i Tammerfors .
När det gäller landsbygdsutveckling , som flera av er tagit upp , bl.a.
Redendo Jiménez , motsvarar riktlinjerna väl de två målsättningar som föredraganden nämner : en stark jordbrukssektor , knuten till ökad konkurrenskraft i landsbygdsområdena , men också bevarande av miljön och landsbygdsarvet i Europa .
Det måste emellertid betonas att de riktlinjer vi talar om endast gäller strukturfonderna , där mål 1 och 2 bl.a. prioriterar diversifiering av landsbygden .
Men när det gäller denna balans på landsbygden får vi heller inte glömma den nya politiken för landsbygdsutveckling , som samfinansieras av Europeiska utvecklings- och garantifonden för jordbruket ( EUGFJ ) garantisektionen , och vars roll är att främja en reformering av det europeiska jordbruket och stödja ett jordbruk med många dimensioner .
Jag skulle på det här stadiet bara vilja säga att jag önskar att det skall införlivas i programplaneringen för landsbygdsområdena inom mål 2 , på samma sätt som EUGFJ : s utvecklingssektion inom mål 1 .
Jag har på den här punkten i vilket fall som helst förstått att man inom utskottet för jordbruk och landsbygdens utveckling är vaksam .
Innan jag slutar skulle jag vilja säga till Savary att i morgon har vi en särskild debatt om konsekvenserna av de stormar som drabbat Frankrike , Österrike och Tyskland framför allt de senaste veckorna , och samtidigt skall vi på nytt , tillsammans med min kollega De Palacio , tala om de lärdomar vi kan dra av oljeutsläppen som också drabbat den franska kusten .
Herr Savary !
Jag avvaktar därför med att ge er min uppfattning , som i stora delar överensstämmer med er egen rekommendation , om vad vi kan göra för att bekämpa detta oljeutsläpp med hjälp av mål 2 .
Jag vill erinra om att kommissionen i morgon skall godkänna kartan över mål 2 för Frankrike , Sverige , Österrike och Luxemburg .
Vi får då ett verktyg för att arbeta bl.a. i en stor del av de områden som drabbats av stormarna .
Det är för övrigt av den anledningen som jag i övermorgon personligen skall resa till två franska departement som allvarligt skadats av stormarna .
Avslutningsvis skulle jag - och jag tackar er herr talman för er förståelse - vilja tacka er , fru föredragande , för det utmärkta arbete som ni och ert utskott utfört , och säga att jag är mycket glad , bortsett från några olikheter när det gäller riktlinjernas roll - vi har talat om det och jag har försökt att klargöra min ståndpunkt - jag är mycket glad över kammarens stöd till kommissionens utarbetande av dessa riktlinjer , som överlämnats till medlemsstaterna för att de skall kunna förbereda sina egna program .
Det kan bara stärka konceptet grundat på ett antal goda tillämpningar efter erfarenheterna från programmen 1994-1999 .
Herr Hatzidakis !
Jag tror det bådar gott för samarbetet mellan våra båda institutioner när nu programplaneringen för 2000-2006 inleds , liksom för goda tillämpningar av samarbete som förstärks av respekten , och det är jag mycket medveten om , för den uppförandekodex som förenar våra två institutioner .
( Applåder ) Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl.12.00.
 
Den sociala och ekonomiska situationen i unionens regioner Nästa punkt på föredragningslistan är debatten om betänkande ( A5-0107 / 1999 ) av Berend för utskottet för regionalpolitik , transport och turism om Sjätte periodiska rapporten om den sociala och ekonomiska situationen i Europeiska unionens regioner [ SEK ( 99 ) 0066 - C5-0120 / 99 - 1999 / 2123 ( COS ) ] . .
( DE ) Herr talman , kommissionär Barnier , mina ärade damer och herrar , kära kolleger !
Den sjätte periodiska rapporten innehåller en omfattande och detaljerad beskrivning av den sociala och ekonomiska situationen i unionens regioner samt deras utvecklingstendenser och bildar , som jag ser det , en solid bas för formuleringen av strukturpolitiska prioriteringar på unionsnivå .
Betänkandet visar att en återhämtningsprocess - mätt i bruttonationalinkomst per capita - har ägt rum och också fortgår i de fattigaste regionerna .
Detta kan till stor del förklaras av strukturfonderna , även om skillnaderna mellan de fattigaste och de rikaste områdena fortfarande är avsevärda .
I och med tillämpningen av de europeiska strukturfonderna har en tillnärmning av levnadsförhållandena skett .
Skillnaderna i den genomsnittliga bruttonationalinkomsten har minskat med 10 procent på tio år .
Särskilt drabbade - givetvis i positiv mening - är de fyra sammanhållningsländerna och även de fem nya tyska förbundsländerna .
Tyvärr har denna utveckling över hela Europa huvudsakligen skett genom en stegring av produktiviteten och endast i liten utsträckning genom sysselsättningstillväxt .
Därför uppmanar vi kommissionen och medlemsländerna att i framtiden ta nödvändig hänsyn även till hur åtgärderna inverkar på sysselsättningen .
Huvuddelen av överföringarna har använts och används för rationaliserings- och moderniseringsinvesteringar för att förbättra arbetsproduktiviteten .
Detta har dock i motsvarande mån dämpat effekterna av den strukturella sysselsättningspolitiken .
Detta är ingen bedömning utan för tillfället ett rent konstaterande .
Betänkandet visar emellertid att de regionala skillnaderna på arbetsmarknaden rentav har fortsatt öka .
I de 25 fattigaste regionerna uppgår arbetslösheten i dag till 24 procent .
För tio år sedan var den fortfarande 4 procent lägre , dvs .
20 procent .
Och i de 25 bästa regionerna , för att nu även nämna detta , har vi i dag en genomsnittlig arbetslöshet på 3,6 procent , för tio år sedan 2,5 procent , alltså en ökning med endast 1,1 procent .
Betänkandet visar tydligt att 50 procent av arbetslösheten är en strukturell arbetslöshet .
Därför , och det är en slutsats som dras i betänkandet , måste kärnan i strukturpolitiken vara främjandet av konkurrenskraften inom näringslivet , stöd åt en näringslivsnära infrastruktur .
Här är ordningsföljden tillika rangordning .
I sammanhanget måste man - vilket bör sägas i direkt anslutning till detta - nämna inte minst åtgärder för att omskola och vidareutbilda arbetskraften .
Vidare måste man i högre grad vara uppmärksam på att stärka företagarpotentialen i de små och medelstora företagen samt att fortsätta utveckla tjänsterna för de små och medelstora företagen .
En annan slutsats i betänkandet är att stödåtgärderna i enlighet med en effektiv stödmedelsinsats måste anpassas enligt ett brett uppdelat medelklass- och existensgrundande stöd .
En mycket viktig punkt , enligt min åsikt .
I resultatet av betänkandet uppmärksammar vi kommissionen på att det rättsliga underlaget för ett samarbete mellan regioner och medlemsländer och kandidatländer måste förbättras samt pekar på det särskilt nödvändiga med en budgetkonsolidering som förutsättning för att den ekonomiska och monetära unionen liksom utvidgningen österut skall kunna lyckas .
Vi uppmanar de medlemsländer som ännu inte har lämnat in en godkänd utvecklingsområdeskarta att göra detta omgående och förväntar oss förstås vidare att kommissionen i ljuset av resultaten från den sjätte periodiska rapporten snabbt granskar regionernas operativa program för den nya stödperioden 2000 till 2006 samt gör allt för att stödperioden också skall kunna dras igång ordentligt och utan förseningar på plats .
Herr talman , herr kommissionär , kära kolleger !
Denna sjätte periodiska rapport om den sociala och ekonomiska situationen i Europeiska unionens regioner innebär ett framsteg i analysen av de regionala uppgifterna och belyser vad som hittills åstadkommits på området , sedan den femte periodiska rapporten kom ut .
Jag anser emellertid att påståendet att de europeiska regionerna genomsnittligt ligger på samma utvecklingsnivå utgör en något stympad bild av situationen , och tyvärr är det ofta vad som återges i pressen och i vissa tal .
Kommissionens rapport sätter till stor del detta påstående i sitt sammanhang , bl.a. när den tar upp den sociala och ekonomiska situationen för vissa regioner inom unionen som ligger mig särskilt varmt om hjärtat : jag tänker på de utomeuropeiska franska departementen och , rent generellt , de yttersta randområdena .
Jag gläds därför åt att utskottet för regionalpolitik antagit ett av mina ändringsförslag som uppmanar kommissionen att avsätta ett eget kapitel i den kommande rapporten om sammanhållningen för de yttersta randområdena , närmare bestämt till att analysera effekten av de åtgärder som inom kort kommer att antas genom tillämpning av den nya artikel 299.2 i Amsterdamfördraget .
Avslutningsvis förefaller det mig som om den sjätte periodiska rapporten innehåller intressanta argument inför ett verkligt projekt för hållbar och rättvis utveckling av det europeiska territoriet , bl.a. när den sammanfattar betydelsen av förhållandet mellan Centraleuropa och de yttersta randområdena .
Även om kommissionen fortfarande tvekar att säga det alltför tydligt visar den periodiska rapporten att vi snarast måste främja en utveckling av gemenskapen med flera olika utvecklingscentrum , via unionens strukturpolitik och inom ramen för de åtgärder som inletts genom SEK ( det europeiska nationalräkenskapssystemet ) .
Herr talman !
Europeiska socialdemokratiska partiets grupp i detta parlament ställer sig bakom det betänkande som Berend just har lagt fram och vi gratulerar upphovsmannen , både till hans fina slutsatser och till hans flexibilitet som har gjort det möjligt för utskottet att införa ändringsförslag från de olika grupperna .
Vi bör ha i åtanke att Europeiska unionens totala konkurrenskraft utgör 81 procent av konkurrenskraften i Förenta Staterna , och att denna siffra endast kan förbättras om den gör det i våra konkurrensdugliga enheter , det vill säga i regionerna , och detta i en tid då den tekniska utvecklingen , internationaliseringen av ekonomin och de problem vi har , utvidgningen och den gemensamma valutan kräver en ökad konkurrenskraft av regionerna , men även av företagen och av den enskilde .
Europeiska kommissionens sjätte rapport innehåller värdefulla slutsatser .
Jag vill sammanfatta två av dessa , som föredraganden redan har tagit upp , en positiv och en negativ sådan .
Den första är att betydande framgångar har uppnåtts vad beträffar den territoriella och sociala sammanhållningen i hela unionens territorium , och att gemenskapens fonder har spelat en viktig , om än ej avgörande roll för att minska de regionala olikheterna .
Den negativa slutsatsen är att de omfattande insatserna har lett till bättre resultat i fråga om utjämningen av BNI och produktiviteten i de europeiska regionerna än i fråga om sysselsättningen .
Därför är det viktigt att den strukturella finansieringen i större utsträckning kopplas till skapandet av arbetstillfällen .
Det , herr kommissionär , är det främsta budordet för den kommande perioden .
Slutligen vill jag , herr talman , uppmana mina kolleger att anta detta betänkande , och i likhet med andra kolleger ber jag kommissionen beakta slutsatserna i den sjätte periodiska rapporten vid utformningen av programmet för åren 2000-2006 .
Herr talman , herr kommissionär , bästa kolleger !
För det första vill jag tacka föredraganden för ett bra arbete och också för att han på ett sakligt sätt beaktat ändringsförslagen under utskottsbehandlingen .
Den sjätte periodiska rapporten lägger grunden för en bedömning av hur unionens regionalpolitiska mål uppnåtts .
Rapporten visar att tillväxten trots alla ansträngningar är ojämn .
Den mycket snabba tillväxten i de centrala delarna av Europa fortsätter .
De starkaste centra växer också hela tiden snabbare än det europeiska genomsnittet , medan utvecklingen i många sydeuropeiska och nordliga regioner går betydligt långsammare .
Nu behövs en djupgående analys av varför regionalpolitiken inte leder till önskat resultat i alla regioner .
Är det byråkratin som är boven eller har man inte i tillräcklig utsträckning tagit hänsyn till skillnaderna mellan regionerna , de långa avstånden , det för kalla eller för varma klimatet , den glesa bebyggelsen och de karga förhållandena ?
På vilket sätt kan unionen möta de utmaningar som den globala utvecklingen medför , så att de svagare utvecklade regionerna kan hänga med i utvecklingen ?
Det är också viktigt att utreda hur unionens utvidgning kommer att påverka strukturfonderna och utvecklingen av unionens randområden .
Medlemsstaterna måste också komma ihåg sitt eget ansvar .
Somliga medlemsstater har brutit mot ökningsprincipen och minskat sina nationella regionala medel när regionalstödet från unionen ökat .
Detta har tärt på regionalpolitikens resultat .
I fortsättningen måste man också fundera på att utveckla indikatorer för att åtgärderna skall kunna riktas in på rätt plats vid rätt tidpunkt .
Man har till exempel inte i tillräcklig utsträckning tagit hänsyn till den okontrollerade migrationen .
Även i detta sammanhang finns det skäl att framhålla de små och medelstora företagens avgörande roll som skapare av sysselsättning och som den regionala utvecklingens motor .
Alldeles speciellt viktigt är det att överföra den nyaste tekniken och ställa know-how till företagens förfogande i de områden där utvecklingen går långsammare .
Vår grupp ställer sig bakom detta betänkande .
Herr talman , herr kommissionär , ärade ledamöter !
Europeiska unionens regionalpolitik har hittills inte lyckats förändra de befintliga skillnaderna i inkomst per capita .
Situationen är allvarlig , vi har alltså i dag i Europeiska unionen en tydlig relation mellan arbetslöshet och fattigdom , vilket visas av det mycket oroande faktumet att arbetslösheten uppgår till i genomsnitt 23,7 procent i de mest drabbade regionerna , regioner som sammanfaller med fattiga regioner , medan arbetslösheten i de 25 områden med minst arbetslöshet , vilka ligger i de rika regionerna , bara uppgår till 4 procent .
Med hänsyn till denna situation bör behovet av åtgärder ämnade att bekämpa den relativa fattigdomen och arbetslösheten klart framgå i det betänkande parlamentet skall godkänna .
Åtgärder som exempelvis en riktig tillämpning av strukturfonderna , vilka ofta används felaktigt , för dessa ändamål , genom en central statlig politik , modernisering av telekommunikation och kommunikationer , särskilt genom att integrera de mindre utvecklade områdena i de transeuropeiska järnvägsnäten med inriktning på år 2007 , respekten för och utvecklingen av jordbrukets och fiskets resurser och förmåga i dessa länder , vilka ofta angrips av Europeiska unionens egen okänsliga politik , samt främjandet av en aktiv sysselsättningspolitik , framför allt för kvinnor och ungdomar .
Bara med en beslutsam tillämpning av denna typ av åtgärder kan man komma över en social och geografisk ojämlikhet som inte är en historisk produkt av oundvikliga misstag , utan tvärtom av en marginalisering och en ekonomisk politik med negativa effekter . )
Herr talman , herr kommissionär !
Berends betänkande följer exakt den strategi som Europeiska kommissionen har definierat genom att frågan om ökad konkurrenskraft ställs i absolut fokus .
Det övergripande målet med strukturfonderna , som till exempel skapandet av fler arbetstillfällen , höjd garanti så att alla bereds samma möjligheter , stabilare villkor för sysselsättning och utveckling , nämns endast i förbigående .
Detta synsätt förefaller mig oberättigat , och jag ber om att större vikt läggs vid dessa punkter i den sjunde periodiska rapporten .
Detta betyder inte att jag inte skulle inse det nödvändiga i att vara konkurrenskraftig , snarare tvärtom i och med att jag själv är företagare i ett mål 1-område , i Brandenburg i förbundsrepubliken Tyskland , och mycket väl känner till de små och medelstora företagens oro och bekymmer .
I mål 1-regionerna är det parallellt med detta absolut nödvändigt med tidsbestämda åtgärder , och då menar jag åtgärder för att skapa nya jobb , särskilda program för att främja förvärvsarbete bland kvinnor och initiativ för att underlätta för den som vill starta eget .
Detta stöds genom lämpliga åtgärder från Europeiska unionens strukturfonder .
Bara genom att stödja företagens konkurrensduglighet kompenserar man aldrig den eftersträvade sammanhållningen mellan ekonomisk och social utveckling , eftersom det helt enkelt saknas grundförutsättningar för en självbärande utveckling i mål 1-regionerna .
Och erfarenheten att den ekonomiska utvecklingen inte själv bidrar till att avskaffa arbetslösheten stöds ju av det faktum att man behöver en ökning av BNP på minst 3 procent för att över huvud taget skapa några nya arbetstillfällen .
Den ensidiga koncentrationen på en ekonomisk politik orienterad efter tillgång , efter efterfrågan kan inte fungera så .
Och driver man en sådan politik måste man satsa mer på utvidgning och mindre på rationalisering .
Man måste absolut länka samman detta med en ekonomisk politik som orienteras efter efterfrågan för att vi alls skall ha en chans att förbättra den sociala situationen i dessa områden .
Situationen skiljer sig markant från region till region .
Det betyder att det krävs en mängd ytterligare åtgärder för att man alls skall kunna åstadkomma något .
Detta vore exempelvis åtgärder för att främja yrkesutbildning , vidareutbildning , för att hjälpa till och slussa tillbaka människor som stötts ut från produktionsprocessen , en flexibel utformning av arbetstid och arbetsformer för att jämka ihop personliga och sociala aspekter på ett avgjort bättre sätt och kanske , återigen , för att främja kvinnors plats i förvärvsarbetet .
Herr talman !
Mina komplimanger till föredraganden för hans ingående betänkande .
Huvudmålsättningen för strukturfonderna är att öka den sociala och ekonomiska sammanhållningen mellan regionerna inom Europeiska unionen .
Genom att stimulera investeringar av olika slag försöker Europeiska unionen att förverkliga en ökning av BNP per capita och en ökning av sysselsättningen .
Av den sjätte periodiska rapporten om regionerna kan man dra den försiktiga slutsatsen att dessa stimulanser inte alltid har den önskade effekten .
Insatserna som syftar till en ökning av BNP per capita i mål 1-områdena resulterar inte alltid i denna ökning .
Det kan inte sägas vara ett tillfredsställande resultat under en period där , framför allt under de senaste åren , ekonomisk framgång varit aktuell .
Såsom föredraganden anger har dessutom effekterna av strukturåtgärderna varit ringa vad sysselsättningen beträffar .
Då är det också på sin plats med en viss återhållsamhet i fråga om gemenskapsstödets effektivitet .
Även konstaterandet att skillnaderna mellan regionerna inom medlemsstaterna ibland rentav ökar väcker allvarliga frågor .
Herr talman !
Det förefaller mig därför vara meningsfullt och nödvändigt att rikta uppmärksamheten , just där det handlar om stimulering av sysselsättningen , såväl på de nationella som på de regionala myndigheterna .
Det är ju de som besitter den största kunskapen om de regioner som faller under deras ansvar .
Genom att låta dem utveckla skräddarsydda planer för de ifrågavarande regionerna och som komplement till detta , om det är nödvändigt , bevilja ekonomiskt stöd kan man uppnå ett bättre resultat .
Och det är ju det som är målet i slutändan .
Därför har jag ingenting att invända mot att kommissionen kommer att överlåta det praktiska utarbetandet och genomförandet av åtgärder till medlemsstaterna och regionerna .
Det är i anslutning till detta möjligen också mer meningsfullt att över huvud taget lägga en större tyngdpunkt på medlemsstaterna med avseende på det ekonomiska stödet till regioner .
Genom att lägga om kriterierna från regionerna till medlemsstaterna förebygger vi en mängd framtida problem .
Slutligen vill jag rikta uppmärksamheten på de central- och östeuropeiska ländernas ställning .
Av betänkandet framgår det att de i allmänhet ligger rejält efter Europeiska unionens länder , i synnerhet på området BNP per capita .
Med tanke på den planerande anslutningen inom överskådlig tid för ett stort antal av dessa länder är det absolut nödvändigt att revidera den nuvarande strukturpolitiken .
Jag vill härmed , efter andras förebild , också uppmana kommissionen att skyndsamt lägga fram förslag till en revidering .
Ärade herr talman , kära kolleger , herr kommissionär !
Efter att noggrant ha studerat föreliggande betänkande måste man tvivelsutan dra slutsatsen att det uppsatta målet med strukturpolitiken har kunnat uppfyllas endast till vissa delar .
Bland annat har klyftorna mellan regionerna snarare ökat än minskat , medlemsstaterna själva registrerar här ett visst närmande .
Likaså har arbetslöshetssiffrorna i de hårdast drabbade regionerna knappast kunnat sänkas , på sina håll har de till och med stigit .
Följaktligen frågar jag mig vad det beror på att anslagen från strukturfonderna inte har använts mer effektivt .
Inte ens kumuleringen av kapitalet från Sammanhållningsfonden och strukturfonderna har varit så framgångsrik i alla regioner som man skulle önska .
Eftersom det nu , över hela Europa , är alla politikers uttalade mål att sänka arbetslösheten måste man ställa en kritisk fråga huruvida den politik som förs är den rätta eller om det är mindre lämpligt att stärka regionernas konkurrensförmåga genom vederbörliga åtgärder såsom ökat stöd åt forskning och utveckling , förbättrad infrastruktur , höjd utbildningsnivå ?
Seriösa strukturreformer och en konkurrensvänligare skatte- och utgiftspolitik är byggstenarna i ett framgångsrikt ekonomiskt säte .
Om vi inte vill låta oss förebrås för att driva en kostnadsintensiv strukturpolitik som inte åstadkommer något varaktigt i sysselsättningsfrågan måste vi analysera hittillsvarande åtgärder .
Unionens strukturpolitik kan betraktas som framgångsrik i och med att man lyckas skapa tillräckligt många arbetstillfällen och arbetslöshetssiffrorna sjunker markant .
Herr talman , herr kommissionär , bästa kolleger !
Jag tackar föredraganden för behandlingen av denna mycket viktiga fråga , för den sociala och ekonomiska situationens utveckling kommer att avgöra hur den europeiska allmänheten bedömer att vi har lyckats i vårt arbete .
Denna fråga , som påverkar människornas vardag , är en nyckelfråga när det gäller Europeiska unionens trovärdighet .
Man måste medge att EU redan har stött utvecklingen i fattiga länder , jag skulle till och med säga att den gjort det på ett storslaget sätt .
Jag minns hur det såg ut i Portugal och i Grekland när jag tävlade där för första gången för tjugofem år sedan .
I detta sammanhang säger nog de som talar franska till EU " coup de chapeau " , dvs. jag lyfter på hatten .
EU är verkligen värd en eloge , men skillnaderna mellan fattiga och rika regioner inom länderna är fortfarande för stora .
Vad blir konsekvensen ?
Folk reagerar genom att rösta med fötterna , genom att ge sig iväg , på jakt efter bröd .
Därför tvingas vi att för samma människor i ett och samma land bygga skolor , sjukhus , hela infrastrukturen om och om igen .
Detta är oerhört dyrt och skapar också mycket stora sociala problem .
De allra flesta skulle dock vilja bo kvar i sin födelsebygd om de fick möjlighet till det , dvs. om det fanns arbete där .
Vi måste ge dem denna möjlighet .
Detta är EU : s och vår moraliska skyldighet .
Som lösning ser jag en klar uppmuntran till företagsamhet .
Med företagsamhet menar jag ingalunda bara att man äger ett företag utan jag menar ett viljemässigt tillstånd .
Jag menar den inställningen att en människa vill gå framåt i sitt liv oavsett om hon är arbetare , företagare eller tjänsteman .
Hur ser ett rättvist samhälle ut ?
Ett samhälle där en människa från enkla förhållanden kan gå framåt i sitt liv för att hennes barn skall få det litet lättare .
På det sättet är det också möjligt att utveckla regionerna i en positiv riktning , för människorna är företagsamma och arbetar om man ger dem möjlighet till det .
Avslutningsvis skulle jag vilja säga att vi i detta fall borde ta lärdom av Amerika där fliten fortfarande står högt i kurs och framgång är ett bevis på kompetens och inte ett föremål för avundsjuka , som ofta är fallet hos oss i Europa .
Herr talman , herr kommissionär , kära kolleger !
Eftersom jag har begränsat med tid skall jag bara ta upp det viktigaste .
Vi kan först och främst konstatera att resultatet av tillväxten inte är rättvist fördelat inom unionen .
Ett exempel är de yttersta randområdena , som fortfarande är hårt drabbade av mycket hög arbetslöshet .
La Réunion har exempelvis en arbetslöshet på 37 procent .
Men det beror inte på konjunkturen utan det är fråga om en strukturmässig arbetslöshet .
Den skapas av det faktum att vi befinner oss långt bort och är en öregion , kort sagt det beror på vår personlighet .
För att bemöta detta innehöll artikel 299.2 i Amsterdamfördraget en princip om särskild och undantagsmässig behandling .
Nu återstår att omsätta denna princip i handling .
Kommissionens dokument som skulle komma i december 1999 har skjutits upp till januari och sedan till februari , och de första kommentarerna gör mig knappast optimistisk .
Jag vänder mig därför högtidligen till rådet och kommissionen .
När det gäller skattefrågor , statligt stöd , strukturfonderna eller att försvara våra traditionella produkter måste vi snarast utarbeta konkreta åtgärder som är både djärva och ambitiösa .
Annars kommer konvergens och sammanhållning tyvärr bara att vara tomma ord , och det finns risk för att den strukturpolitik som bedrivs i våra regioner slutar med ett misslyckande trots att det handlar om så stora belopp . .
( FR ) Herr talman !
Jag skulle i min tur , liksom alla andra talare , vilja tacka herr Berend och lyckönska honom till ett utmärkt arbete .
Liksom när det gäller det tidigare betänkandet är analysen mycket kompetent och exakt , och rekommendationerna , liksom era egna kommentarer mina damer och herrar , kommer att vara till nytta för kommissionen i allmänhet , och för kommissionären med ansvar för regionalpolitik i synnerhet , när vi skall inleda programplaneringen i fråga om anslagen för 2000-2006 .
Jag skulle i min tur vilja göra några kommentarer , till att börja med om er bedömning , herr föredragande , av denna sjätte periodiska rapport .
Ni betonade dess kvalitet och ni skrev till och med , om jag inte misstar mig , att i jämförelse med de tidigare var den betydligt bättre .
Jag vill för kommissionens räkning och för min företrädares , Wulf-Mathies räkning , säga att vi var mycket glada över denna bedömning från kammaren och er .
Kommissionen har verkligen ansträngt sig , herr Berend , för att denna sjätte periodiska rapport skulle göra det möjligt att konstatera en insats , ett kvalitativt steg framåt , i den analys vi föreslår er .
Jag tänker särskilt på innehållet i kapitel 2.1 i rapporten , där kommissionen på ett fördjupat sätt granskat de ekonomiska definitionerna av den regionala konkurrenskraften och försökt analysera hur denna konkurrenskraft kan stödjas , förbättras och påverkas av faktorer som vissa av er , Markov nyss eller Raschhofer , kraftigt betonat .
Jag tänker på teknisk forskning och utveckling , infrastrukturens tilldelning och kvalitet , de mänskliga resursernas potential , de små och medelstora företagen och direktinvesteringar från utlandet .
Så långt kvaliteten .
Herr föredragande !
Jag vill inte nu lägga alltför mycket tid på detaljer om min uppfattning inom olika allmänna punkter där kammaren redan är överens med oss .
Jag skall bara kort nämna dem : den första gäller betydelsen av rapportens slutsatser för att utarbeta prioriteringar för den nya regionalpolitiken , särskilt för förhandlingar om programplaneringsdokument med medlemsstaterna .
Den andra punkten , partnerskapen , som flera av er betonat , handlar om rollen för de lokala och regionala myndigheterna , den privata sektorn , arbetsmarknadens parter samt föreningarna och lokala grupper .
När det gäller problemet med partnerskap kommer jag att mycket noggrant se till att bestämmelserna i den allmänna förordningen om strukturfonderna tillämpas korrekt .
Den tredje punkten gäller behovet av att öka sysselsättningens andel av tillväxten , även om jag mycket väl vet , och van Dam sade det också nyss , att det i första hand är medlemsstaterna som är ansvariga , och att man , när man talar om medlemsstaternas ansvar , liksom om nyttan och effektiviteten av denna regionalpolitik , också måste titta på var vi befinner oss .
Fruteau förklarade nyss att resultatet av tillväxten är orättvist fördelat .
Herr parlamentsledamot !
Det måste ändå finnas en tillväxt och vi kan inte befinna oss i en period av fullständig stagnation eller tillbakagång , vilket förekommit tidigare .
Tillväxt och fattigdom gäller inte alla , kanske ni hävdar .
Jag håller med er .
När tillväxt är ett faktum måste den vara bättre fördelad , men det som är ännu svårare och drabbar de regioner som är avlägset belägna , de yttersta randområdena eller öregionerna ännu allvarligare , är avsaknaden av tillväxt som varit kännetecknade för de två senaste decennierna .
Den fjärde punkt som Hedkvist Petersen nyss betonade är främjandet av en politik för lika möjligheter för män och kvinnor .
Den femte punkten gäller de små och medelstora företagens betydelse och roll , vilket Vatanen starkt betonade nyss .
Slutligen har vi den positiva effekten av strukturfondernas förvaltningssystem på de nationella myndigheterna , tjänstemännens motivation när de förvaltar dessa fonder , även om det ibland är komplicerat , och betydelsen av att på nytt förbättra förfarandet för kommissionens utvärdering , uppföljning och kontroll .
Jag vill i det sammanhanget informera Europaparlamentet om min avsikt att i mitten av år 2000 arrangera ett seminarium med nationella och regionala myndigheter om denna fråga om utvärdering av förfarandena för utbyte av goda tillämpningar när det gäller att förvalta strukturfonderna .
Jag skulle vilja ta upp några specifika punkter .
Herr Berend !
Ni ville att zonindelningen skulle genomföras snabbt .
Vi har avslutat den .
I morgon kommer fyra nya länder att vara föremål för kommissionens beslut och mycket snabbt , hoppas jag , är det Italiens tur .
Ni kommer alltså att bli nöjd på den punkten eftersom alla länder som berörs av mål 2 blir indelade i zoner .
När det gäller den informella ekonomin som ni tar upp i ert betänkande , vet jag naturligtvis att analys och framtagning av statistik på detta område är beroende av uppgifternas tillförlitlighet och såsom Cocilovo också sade föreligger det ett tillförlitlighetsproblem när det gäller dessa uppgifter .
I viss utsträckning beaktas de på nytt i statistiken över BNI och undersökningar om arbetskraften och i vilket fall som helst vill jag betona de ansträngningar Eurostat gör och kommer att göra för att förbättra statistikens kvalitet .
Herr Berend !
Liksom Aparicio Sánchez tog ni upp avsaknaden av reformer på fiskeområdet .
På denna punkt , som personligen intresserar mig , vill jag erinra om att denna sektor är liten - vilket inte betyder att den är betydelselös - och att den är koncentrerad till ett mycket litet antal regioner , och det gör det inte lättare att analysera den inom en regional ram .
Denna typ av sektorsanalys faller mer under generaldirektoratet för fiske , under min kollega Fischlers ledning .
Jag vill ändå försäkra er om att kommissionen kommer att försöka införliva en sådan analys i den andra rapporten om sammanhållningen , som sannolikt bättre kommer att motsvara denna oro .
Flera av er har nämnt punkter som bör ingå i denna andra rapport om sammanhållningen , och föredraganden tog upp några av dessa .
Jag vill till att börja med försäkra er om att sammanslagningen av de periodiska rapporterna och rapporten om sammanhållningen inte på något sätt kommer att innebära att information går förlorad eller att intresset minskar för innehållet i rapporten om sammanhållning som för mig , herr föredragande , är ett mycket viktigt instrument , inte bara för att man redogör för vad som gjorts och gör det på ett öppet och noggrant sätt , eller för att man granskar eller utvärderar kommande riktlinjer , utan också för att skapa en allmän debatt med medborgarna och även med er som folkvalda om denna regionalpolitik och om det som en dag skulle kunna bli en europeisk politik för fysisk planering .
Jag har i vilket fall som helst noterat att ni önskar införliva följande punkter i rapporten : definition , insamling och analys av beståndsdelar som är representativa för regionen och för alla länder i Central- och Östeuropa , ett kapitel om de yttersta randområdena och öregionerna som flera av er tagit upp , särskilt Sudre och Fruteau , analys av regionernas konkurrenskraft i länderna i Central- och Östeuropa - det blir den stora utmaningen för oss , för er , för kommissionen , under de kommande åren , och slutligen de gränsöverskridande aspekterna .
På alla dessa punkter skall jag försöka följa era rekommendationer .
Jag skulle slutligen vilja ta upp några politiska slutsatser som ni för övrigt känner till , men där jag ändå skulle vilja erinra om de viktigaste beståndsdelarna .
Mina damer och herrar !
Avsevärda framsteg har gjorts för att uppnå en verklig konvergens , bl.a. för de fyra sammanhållningsländerna , men också , herr Pohjamo , det säger jag ärligt , för regionerna inom mål 2 som tagit igen viss försening i sin utveckling , bl.a. när det gäller infrastruktur .
Det är den första politiska punkten .
Den andra politiska punkten , strukturfonderna , har lämnat och kommer att lämna ett betydande bidrag till denna tillnärmningsprocess .
Alla makroekonomiska modeller som vi arbetar efter visar för det senaste decenniet att mer än en tredjedel av den konvergens som uppnåtts i regioner med försenad utveckling inte skulle ha ägt rum om det inte vore för strukturfonderna .
Jag har emellertid noterat , när det gäller framför allt de yttersta randområdena , fru Sudre , herr Fruteau , och även herr Nogueira Román , att ni konstaterar att mycket fortfarande återstår att göra - och det är min tredje punkt - när det gäller att öka sysselsättningen , förbättra kampen mot social utslagning , som är särskilt allvarlig och oacceptabel i många av våra regioner samt underlätta för kvinnor och ungdomar att komma in på arbetsmarknaden .
Den fjärde politiska punkten gäller unionens utvidgning , som är det stora politiska och humanistiska projektet för våra institutioner under de kommande åren , och även en stor utmaning för Europas sammanhållningspolitik , en punkt som van Dam betonade .
Jag tror att redan i Berlin och i de finansiella instrument som ställs till vårt förfogande kan man ana det som skulle kunna bli en sammanhållningspolitik för de första nya länder som skall bli medlemmar .
Jag tänker särskilt på ISPA-instrumentet som det är mitt ansvar att genomföra under de kommande veckorna .
Mina damer och herrar !
Som ni ser har vår nya programplanering knappt inletts och vi har redan en gemensam diskussion om effekten av unionens utvidgning på vår strukturpolitik .
Denna sjätte periodiska rapport som ni , herr Berend , totalt sett uttalat er positivt om utgör för oss , för mig , en bra bas för diskussionerna .
Jag skulle därför vilja tacka er mycket uppriktigt för ert bidrag till diskussionerna som vi inlett för de kommande riktlinjerna , liksom för den goda tillämpningen av riktlinjerna för perioden 2000-2006 .
Tack så mycket , herr kommissionär .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
( Sammanträdet avslutades kl .
20.25 . )
