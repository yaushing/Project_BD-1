 
Återupptagande av sessionen Jag förklarar Europaparlamentets session återupptagen efter avbrottet torsdagen den 3 februari 2000 .
 
Justering av protokollet från föregående sammanträde Protokollet från sammanträdet torsdagen den 3 februari har delats ut .
Finns det några synpunkter ?
Jag förstår av er reaktion att många av parlamentsledamöterna inte fått protokollet , och det är självklart att ni inte kan justera ett protokoll som ni inte har fått .
Jag föreslår därför att vi justerar det i morgon förmiddag , eftersom ni uppenbarligen inte fått det och det ber jag om ursäkt för .
Justeringen av protokollet skjuts alltså upp .
Fru talman !
Rörande en ordningsfråga .
I förmiddags rapporterade BBC att en brittisk ledamot av Europaparlamentet , som innehar en hög position inom sin delegation , fortsätter att erbjuda strategisk rådgivning till privata klienter , men inte meddelar i intresseregistret vilka dessa klienter är .
Europas medborgare har rätt att förvänta sig att deras företrädare håller isär sitt privata vinstintresse från det allmännas bästa , men de kan bara vara säkra på att detta görs i varje enskilt fall om informationen både är tillgänglig för allmänheten och lätt åtkomlig .
Fru talman !
Eftersom dessa frågor för närvarande diskuteras i kvestorskollegiet , får jag be er att använda ert inflytande både för att se till att intresseregistret uppdateras och ändras för att omfatta fall av denna typ och , framför allt , för att se till att registret inte bara är tillgängligt för inspektion av denna kammare , utan att det också offentliggörs på Internet ?
Tack , herr Davies .
Jag skall titta på frågan med kvestorerna .
Fru talman !
Rörande en ordningsfråga .
Eftersom detta är årtusendets första Alla hjärtans dag , hoppas jag att ni kan hålla med mig om att det skulle vara lämpligt om denna kammare markerade denna dag genom att på ett bestämt sätt åta sig att komma till rätta med hjärtsjukdomarna , vilka orsakar de flesta dödsfallen i Europeiska unionen .
Jag vill uppmana ledamöterna att underteckna det åtagande som gjordes i dag vid the Winning Hearts Conference , att alla barn som föds under det nya årtusendet skall ha rätt att leva i åtminstone 65 år utan att behöva lida av kardiovaskulära sjukdomar som är möjliga att undvika .
Jag önskar er en trevlig Alla hjärtans dag !
( Applåder ) Fru talman !
Jag uttalar mig enligt artikel 9 i denna kammares arbetsordning och åsyftar samma fråga som togs upp av Davies om de mycket allvarliga anklagelserna som uttalades på BBC i förmiddags .
Jag skulle välkomna en försäkran från er att ni kommer att beställa en undersökning för att se till att de två ledamöter som nämndes i denna specifika BBC-intervju inte driver sina företag från detta parlament eller från parlamentets lokaler , eftersom detta i sanning skulle vara mycket allvarligt .
Under årens lopp har de brittiska konservativas dubbelmoral gjort att det brittiska underhuset fått ett dåligt rykte , och det finns en verklig fara att ett sådant uppförande skulle få liknande effekter för detta parlament .
Tack , herr Murphy .
Som jag sade till Davies skall jag redan i kväll titta på frågan tillsammans med kvestorerna .
Fru talman !
Rörande en ordningsfråga .
Jag har redan skrivit till er vid ett flertal tillfällen om hur ordningsfrågor tas upp i kammaren .
Jag undrar vilken ordningsfråga Davies tog upp .
Varför nämnde han inte att en av hans egna liberala kolleger också bedriver rådgivningsverksamhet som håller på att undersökas av BBC ?
Skall denna kammare låta sin föredragningslista bestämmas av plumpa rapporter om ett program som grundar sina nyhetsinslag på lögner , eller skall den utföra ett seriöst arbete och ta itu med de utmaningar som Europa står inför ?
Kära kolleger !
Det är självklart att kvestorerna som skall granska frågan inte enbart kommer att förlita sig på information som hörts i radion .
De kommer att gå igenom detta mycket noggrant .
Fru talman !
Jag tror att jag gör mig till tolk för ett stort antal kolleger i de flesta politiska grupperna när jag säger att det budskap som kommissionens ordförande framförde för en vecka sedan till den nya österrikiska förbundskanslern skapade obehag .
Var det verkligen nödvändigt att säga , jag citerar : " mina varmaste lyckönskningar följer er " , eller " jag betvivlar inte att ni kommer att fortsätta era föregångares engagemang när det gäller frihet och demokrati samt respekt för de mänskliga rättigheterna och grundläggande friheterna " , eller " jag ser fram emot ett fruktbart och konstruktivt samarbete " ?
Fru talman !
Jag skulle vilja att Prodi i morgon berättar för oss vad han ville eller inte ville ge för betydelse åt sitt uttalande så att ingen , absolut ingen , kan utnyttja detta minst sagt bisarra och olyckliga budskap , även mot Prodis vilja , för att bidra till att banalisera den farliga politiska process som äger rum i Österrike .
Tack , herr Wurtz .
Kära kolleger !
Jag ber er att inte inleda någon debatt , det handlade om ett förslag som rör förfaranden .
Jag vill erinra er om , herr Wurtz , att vi i morgon träffar Prodi som kommer att uttala sig om kommissionens program .
Ni har naturligtvis full frihet att i era inlägg efter uttalandet fråga ut honom , på samma sätt som Prodi har fullständig frihet att svara er .
Jag föreslår att vi definitivt klargör denna fråga då , om ni och Prodi vill det .
Fru talman !
Jag är mycket ledsen över att jag återigen måste besvära er med en punkt som jag redan tagit upp här två gånger tidigare .
Jag har redan talat om för er ett antal gånger att vi för de nederländska kollegernas räkning gärna skulle vilja ha en nederländsk TV-kanal .
Det finns nu 28 kanaler här i parlamentet , därav två grekiska , en portugisisk , en finsk och en belgisk , men fortfarande ingen nederländsk , däremot sju engelska , sex tyska och sex franska .
Redan i september fick jag löfte om att det skulle finnas en nederländsk kanal i januari .
Det är nu februari , och det finns fortfarande ingen .
Jag skulle därför återigen vilja be er att vidta åtgärder för detta .
Jag undrar vilken medeltida byråkrati det är som förhindrar att en nederländsk kanal överförs via satellit .
Fru Plooij-van Gorsel !
Jag är också besviken , eftersom jag själv var övertygad om att frågan hade lösts för länge sedan .
Jag har noterat era budskap i frågan och jag tror att Banotti har ett svar till er .
Jag skall därför , om ni tillåter , lämna ordet till Banotti så att hon kan svara er i form av ett förslag som rör förfaranden .
Fru talman !
Som min kära vän Elly vet , kommer jag att göra allt för att se till att hon och mina nederländska kolleger blir nöjda .
Jag kan i egenskap av kvestor med ansvar för denna fråga försäkra er om att vi haft tekniska diskussioner om de olika kanalerna på TV och radio , och jag har redan börjat skicka brev till kolleger i detta ärende .
Om det nu kan lugna henne , har inte irländarna heller fått sin kanal ännu .
Det verkar finnas svårartade tekniska problem , men vi arbetar verkligen på det .
Tack för att jag fick möjlighet att reda ut detta .
Jag är inte säker på att våra nederländska kolleger känner sig lugnade , eftersom våra irländska kolleger inte heller kan få in någon inhemsk kanal .
Jag tror att vi måste titta på vad som kan göras så att alla kolleger kan se sin kanal .
Tack , fru Banotti , och övriga kvestorer , för era ansträngningar i ärendet .
Fru talman !
Jag ville säga till herr Wurtz att kommissionens doktrin inte är Bresjnevs doktrin om begränsad suveränitet och att vi inte , till dess att motsatsen bevisats , befinner oss inom ramen för artikel 6 och 7 .
Österrike har därför fullständig rättighet att bilda en regering och kommissionens ordförande har fullständig rättighet , och till och med skyldighet , att framföra sina lyckönskningar till Österrike .
Wurtz kanske borde erinra sig att det inte var så länge sedan som kolleger i hans parti , franska kommunistiska borgmästare , skickade ut bulldozrar mot invandrarförläggningar i Frankrike .
 
Arbetsplan Nästa punkt på föredragningslistan är fastställande av arbetsplanen .
Det slutgiltiga förslaget till föredragningslista som utarbetats av talmanskonferensen i enlighet med artikel 110 i arbetsordningen har delats ut. a ) Sammanträdet den 14 till 18 februari 2000 i Strasbourg Beträffande onsdagen : Talmannen .
Med tanke på att rådet inte kan vara närvarande onsdag kväll har flera grupper - Europeiska folkpartiet , Europeiska socialdemokratiska partiet , de liberala , De gröna och den enade vänstern - begärt att vi i en gemensam diskussion skall behandla rådets uttalande om den cypriotiska frågan och Broks betänkande om föranslutningsstrategin för Cypern och Malta och flytta fram dessa punkter , liksom Swobodas betänkande i föredragningslistan .
Det skulle alltså innebära att vi på onsdagen har rådets två uttalanden om sammanhållningen mellan unionens politik och utvecklingspolitiken och om FN : s session om " Mänskliga rättigheter " , följt av den gemensamma diskussionen om Cypern och sedan om betänkandena från Swoboda , Frassoni och Knörr Borràs , samt rapporten från Corrie .
Vem vill lägga fram denna begäran i dessa gruppers namn ?
Då ingen begärt ordet låter jag alltså begäran gå till omröstning .
( Parlamentet biföll begäran . ) Beträffande torsdagen : Talmannen .
När det gäller aktuella och brådskande frågor av större vikt har jag mottagit flera önskemål om ändringar .
När det gäller mänskliga rättigheter har jag mottagit två önskemål om tillägg : ett från den liberala gruppen om en underpunkt med beteckningen " Kambodja " och ett från Gruppen De gröna om en underpunkt med beteckningen " Pinochet " .
Som ni vet kan punkten " Mänskliga rättigheter " inte omfatta fler än fem frågor .
Förteckningen i det slutgiltiga förslaget till föredragningslista omfattar nu fyra frågor och vi kan därför bara lägga till ytterligare en .
Vem vill lägga fram begäran om en underpunkt om Kambodja för den liberala gruppens räkning ?
Fru talman !
För den liberala gruppen är det av stor vikt att en diskussion om situationen i Kambodja äger rum , och att det sker just nu .
Inte bara på grund av brevet som Förenta nationernas generalsekreterare , Kofi Annan , skrivit till Kambodjas regering för att den någon gång skall vida åtgärder för en särskild tribunal i syfte att ställa röda khmerernas ledare till svars , utan också för att Hun Sens regim , som uppenbarligen inte är nöjd med mordförsöken på oppositionsledaren Sam Raninsy , nu har kommit på att man kanske kunde upphäva hans parlamentariska immunitet för att han helt enkelt skall kunna ställas inför rätta .
Världssamfundet har krävt att de skyldiga skall ställas till svars för det som sker i Kambodja .
När allt kommer omkring var det vi som godkände valet i Kambodja , vilket måste betecknas som ett av de största fiaskona på området valobservation .
Det var bara parlamentet som kom ur detta med ett visst anseende i behåll .
Jag tror att vi från parlamentets sida måste ta vårt ansvar även den här gången och göra ett uttalande om situationen i Kambodja .
( Parlamentet biföll begäran . )
Talmannen .
Underpunkten Kambodja läggs alltså till under punkten " Mänskliga rättigheter " , vilket gör att begäran om en underpunkt rörande Pinochet inte kan bifallas .
Jag har också mottagit önskemål om att lägga till nya punkter i den aktuella och brådskande debatten om frågor av större vikt .
Det handlar alltså inte längre om att lägga till frågor under rubriken " Mänskliga rättigheter " , utan att lägga till nya punkter .
Jag har mottagit tre önskemål : en första begäran från den enade vänstern om att lägga till en punkt " Moratorium om dödsstraff i Förenta staterna och fallet med Betty Beets " , en andra begäran från den liberala gruppen om att lägga till en ny punkt med beteckningen " Pinochet " , och en tredje begäran från Gruppen De gröna om att lägga till en ny punkt " Katastrofer : Donaus miljö " .
Med tanke på den tid vi förfogar över , och eftersom vi som ni vet har ett uttalande från kommissionen om omstrukturering av företag , och den nuvarande förteckningen omfattar två punkter , kan vi alltså lägga till ytterligare två .
Jag skall först ta begäran från gruppen den enade vänstern .
( Parlamentet avslog begäran . )
Talmannen .
Vi går nu vidare till begäran från den liberala gruppen .
Finns det någon som vill uttala sig för den ?
Fru talman !
Det är påfallande att Europaparlamentet hittills inte har tagit ställning i fråga om det eventuella frisläppandet av Pinochet trots de internationella häktningsorder som redan utfärdats .
Med tanke på att den belgiska regeringens överklagande gillades förra veckan och med tanke på att beslutet i huvudsak ännu inte är fattat är det viktigt att parlamentet äntligen ger en ordentlig signal , en signal som borde innehålla att ingen kan undkomma en rättvis rättegång .
Det är otänkbart att Europaparlamentet , som med rätta ägnar så mycket uppmärksamhet åt respekten för de mänskliga rättigheterna , inte skulle göra något tydligt uttalande i detta fall .
Fru talman !
Detta är en fråga som är alldeles för allvarlig för att i nuläget behandlas som ett brådskande ärende .
För det första har Europaparlamentet redan uttalat sig om general Pinochet , men förutom det måste vi nu påminna oss vissa saker .
Den första är att detta är ett ärende som är sub iudice i flera europeiska länder , och jag påminner kollegerna om att det ännu inte existerar ett europeiskt straffrättsligt område och inte heller ett europeiskt rättsområde .
Vi är för den internationella brottmålsdomstolen , men den finns inte ännu .
För det andra finns det för närvarande en demokratiskt vald regering i Chile , under ledning av Ricardo Núñez , vars första uttalande varit att alla som begått brott av detta slag skall ställas inför rätta .
Och jag påminner mig att den chilenska rättvisan , som är oberoende , för närvarande går igenom 60 stämningsansökningar mot general Pinochet och hans brott mot mänskligheten .
Jag anser att frågan är så viktig att vi bör följa den , men inte att vi skall lösa den med hjälp av förfarandet för brådskande ärenden .
Vi är för att rättvisa skipas i denna frågan , men vi tror inte att det här är det lämpligaste sättet .
( Parlamentet avslog begäran . )
Talmannen .
Vi kommer nu till den tredje begäran som är " Miljökatastroferna i Donaus vatten " , en begäran från Gruppen De gröna .
Finns det någon ledamot som vill lägga fram denna begäran ?
Fru talman , kära kolleger !
Det som hänt i en av Donaus bifloder anses av många specialister som en olycka med samma allvarliga inverkan på miljön som Tjernobylkatastrofen .
Det drabbar inte bara Rumänien , utan också Jugoslavien , det drabbar faktiskt hela Donaudalen .
Vi anser att frågan är tillräckligt allvarlig för att kommissionen snabbt skall reagera på denna situation , och jag anser att parlamentet bör uttala sig och rösta för en resolution i frågan .
( Applåder ) ( Parlamentet biföll begäran . )
Talmannen .
När det gäller torsdagen har PPE-gruppen också begärt att Cederschiölds betänkande om förstärkning av det straffrättsliga skyddet mot förfalskning i samband med införandet av euron skall tas upp som sista punkt på onsdagen .
Finns det någon kollega som önskar uttala sig för PPE-gruppen och lägga fram denna begäran ?
Fru talman !
Jag vill bara be kammaren att stödja detta förslag , eftersom det har varit väldigt många omflyttningar i denna föredragningslista .
Det är ett ganska kort ärende , men det är extremt viktigt att det passerar parlamentet nu , och att det inte blir några förseningar .
Det handlar nämligen om förfalskningar av euron , vilket är ett ärende som är väldigt brådskande .
Vi har försökt driva igenom detta .
Jag vore därför väldigt tacksam om kammaren skulle kunna stödja detta förslag .
( Parlamentet biföll begäran . )
Beträffande fredagen : Talmannen .
När det gäller fredagen har vi på förmiddagen en muntlig fråga om posttjänster och Europeiska socialdemokratiska partiets grupp begär att resolutionsförslagen skall gå till omröstning direkt efter debatten och inte i Bryssel , såsom föreslagits i det slutgiltiga förslaget till föredragningslista .
Vill någon kollega yttra sig för PSE-gruppen och lägga fram denna begäran ?
Fru talman !
Jag ber min vän Enrique Barón om ursäkt , men jag skulle vilja uttala mig emot detta förslag .
Jag är till och med förvånad över att det dyker upp , eftersom vi hade kommit överens om detta efter diskussion i talmanskonferensen .
Fru talman !
Jag tror att ert förslag att dela upp det hela med debatt på fredag och omröstning senare är klokt .
Skälet är följande : frågan berör inte mindre än 1 800 000 löntagare inom Europeiska unionen .
Vi har ett direktiv .
Det är inte gammalt , det härrör från 1997 .
Att inför ett nytt direktiv besluta om den framtida inriktningen i all hast , utan att ha tid att rådfråga fackföreningarna eller diskutera med samtliga parter på arbetsmarknaden , tycker jag strider mot den anda som vi vill ingjuta i debatten om frågor som direkt berör arbetsmarknadens parter .
Jag är alltså för att vi behåller den ursprungliga uppdelningen : debatt på fredag , omröstning senare .
Fru talman !
Det är tydligen så att jag är skyldig Wurtz en förklaring , och jag skall ge hela parlamentet den .
Vi hade nått denna principöverenskommelse i talmanskonferensen .
Jag visste inte då att kommissionär Bolkestein skulle komma nästa vecka för att tala om denna fråga i utskottet för regionalpolitik , transport , och turism .
I min grupp har vi diskuterat frågan och , med beaktande av det nuvarande läget för hela integrationsprocessen av marknaden och avregleringen av en så känslig fråga , anser vi att det är lämpligt att parlamentet gör ett första uttalande , oberoende av vad det gör i framtiden , så att kommissionär Bolkestein kan notera detta och för att ge en inriktning till debatten nästa vecka .
Fru talman !
Jag vill helt enkelt be kollegan Wurtz att läsa igenom vad det här handlar om .
Det är inte fråga om någon innehållslig kontrovers utan endast om frågesatsen : När skall kommissionen , efter att nu ha haft ett och ett halvt år på sig , äntligen vara i stånd att lägga fram direktivet ?
Vad vi vill med resolutionen är bara att de utsatta tiderna skall hållas , och då är det viktigt att vi agerar så snabbt som möjligt .
Därför vill jag stödja socialdemokraternas förslag att genomföra omröstningen på fredag .
( Parlamentet biföll begäran . )
Fru talman !
Cederschiöldbetänkandet avfördes ju från torsdagens föredragningslista .
Därmed torde vi få litet tid över på torsdag .
Eftersom vi , med hänsyn till det stora antal frågor som skall avhandlas på en och en halv timme , ju har mycket knappt om tid för de brådskande ärendena vill jag bara fråga sessionstjänsten om man inte kan undersöka huruvida vi kan få en halvtimme extra för de brådskande ärendena för att få talartiden att räcka .
Det förefaller mig över huvud taget som om fördelningen av sessionstiden de senaste veckorna har varit mycket kaotisk .
Det rådde stor tidspress under talartiderna , men så plötsligt hade vi en till en och en halv timme över förra torsdagen , då inget ämne fanns upptaget på föredragningslistan och vi blev tvungna att vänta på omröstningen .
På fredag i denna vecka har vi ett en fråga .
Det är faktiskt absurt .
Jag vill verkligen be om en granskning av hur ekonomiskt sessionerna planeras .
Det är fullständigt möjligt : låt oss därför se om vi kan förlänga tiden för de brådskande frågorna med en halvtimme , eftersom Cederschiölds betänkande utgår .
Det är vad det handlar om , och enbart detta .
Fru talman !
Jag skulle vilja göra ett inlägg om en punkt på föredragningslistan för onsdagen , som ni inte tagit upp .
Jag förstår att det inte är en polemisk fråga att uttalandet om 50-årsdagen av Genèvekonventionerna inte innefattas i rådets uttalande om nästa möte i Förenta nationernas kommitté för mänskliga rättigheter och att detta uttalande , för att utformas på ett ädelt och högtidligt sätt överlämnats till plenum i mars .
Jag förstår att det finns en överenskommelse om detta .
Fru talman !
Under denna eftermiddag i denna kammare har det hänvisats till en rad rapporter på BBC : s program Today denna förmiddag , i vilket man hävdade att vissa av mina kolleger drev personliga lobbyföretag eller på något sätt missbrukade sin ställning som ledamöter av denna kammare .
Detta är allvarliga anklagelser .
De är fullständigt osanna , ondskefulla , politiskt färgade och de uttalades trots vetskapen om att de var osanna .
Vi skall vidta rättsliga åtgärder .
Mina kollegers intresseregister är fullständiga .
Om vi får vetskap om att någon ledamot av denna kammare eller dennes medarbetare samarbetat med BBC i denna röra kommer vi att avslöja dem , vilket drar skam över denna kammare .
Det stämmer , vi är helt överens. b ) Sammanträdena den 1 och 2 mars 2000 i Bryssel
 
Hållbar stadsutveckling - Landsbygdens utveckling - Equal-initiativet Nästa punkt på föredragningslistan är gemensam diskussion om följande fyra betänkanden : betänkande ( A5-0026 / 2000 ) av McCarthy för utskottet för regionalpolitik , transport och turism om meddelandet från kommissionen till medlemsstaterna om fastställande av riktlinjer för ett gemenskapsinitiativ för ekonomisk och social förnyelse av städer och förorter som befinner sig på tillbakagång för att främja hållbar stadsutveckling ( Urban ) ( KOM ( 1999 ) 477 - C5-0242 / 99 - 1999 / 2177 ( COS ) ) ; betänkande ( A5-0028 / 2000 ) av Decourrière för utskottet för regionalpolitik , transport och turism om kommissionens meddelande till medlemsstaterna med riktlinjer för ett gemenskapsinitiativ som rör transeuropeiskt samarbete och syftar till en harmonisk och balanserad utveckling av det europeiska området ( Interreg ) ( KOM ( 1999 ) 479 - C5-0243 / 99 - 1999 / 2178 ( COS ) ) ; rapport ( A5-0024 / 2000 ) av Procacci för utskottet för jordbruk och landsbygdens utveckling om förslaget till kommissionens meddelande till medlemsstaterna om fastställande av riktlinjer för gemenskapsinitiativet för landsbygdens utveckling ( Leader + ) ( KOM ( 1999 ) 475 - C5-0259 / 99 - 1999 / 2185 ( COS ) ) ; betänkande ( A5-0034 / 2000 ) av Stenzel för utskottet för sysselsättning och socialfrågor om utkastet till meddelande till medlemsstaterna om fastställande av riktlinjer för program inom ramen för gemenskapsinitiativet Equal för vilka medlemsstaterna uppmanas lämna in förslag till stöd ( KOM ( 1999 ) 476 - C5-0260 / 99 - 1999 / 2186 ( COS ) ) .
Eftersom McCarthy är litet försenad p.g.a. sitt flyg föreslår jag att vi först lyssnar till Decourrière . .
( FR ) Fru talman , kära kolleger , herrar kommissionärer och ledamöter av utskottet för regionalpolitik , transport och turism !
Jag har fått i uppdrag att upprätta Europaparlamentets betänkande om programmet för gemenskapsinitiativet Interreg III .
När frågan överlämnades till utskottet granskade vi över 100 ändringsförslag och hittills har 17 ändringsförslag på nytt lämnats in , vissa av dem har redan lagts fram för kommissionen .
Innan vi diskuterar innehållet i den resolution som jag lägger fram skulle jag vilja tala om vilka beståndsdelar jag beaktat och använt som riktlinjer för mitt arbete som föredragande .
Till att börja med vill jag erinra om den roll som gemenskapsinitiativet Interreg har , som grundades på principen om gränsöverskridande och innovation .
Programmet är en drivkraft när det gäller utveckling och den europeiska dimensionen .
Interreg är ett av de fyra gemenskapsinitiativ som planeras för perioden 2000-2006 och kommer att förfoga över det största totalanslaget , nämligen 4,875 miljarder euro , jämfört med 3,604 miljarder för närvarande .
Initiativet Interreg inrättades 1990 och bygger på strävan att förbereda de europeiska regionerna för ett Europa utan gränser , inom ramen för den stora inre marknadens genomförande .
Vid reformen av strukturformerna 1994 och 1996 införlivades nya områden i gemenskapsprogrammet Interreg , vilka bidrog till att utveckla transeuropeiska nät för transport och energidistribution .
Dessa program har främjat gränsöverskridande samarbete , liksom samarbete mellan länder och regioner inom Europeiska unionen , genom att främja en balanserad utveckling av gemenskapsområdet .
Programmet Interreg III är en fortsättning av detta arbete och Europeiska kommissionen överlämnar i dag riktlinjerna för detta till oss , i enlighet med bestämmelserna i rådets förordning ( EG ) nr 1260 från 1999 om allmänna bestämmelser för strukturfonderna .
Programmet är uppdelat i tre områden : område A gäller det gränsöverskridande samarbetet mellan territoriella myndigheter och gränsregioner inom och utanför Europeiska unionen , utifrån gemensamma utvecklingsstrategier och där genomförandet faller under medlemsstaterna och de lokala och regionala myndigheterna , område B gäller samarbete mellan länder och mellan nationella , regionala och lokala myndigheter i flera medlemsstater eller kandidatländer , inom områden som fysisk planering , transport- och miljönätverk .
Genomförandet av detta område är medlemsstaternas och de nationella myndigheternas ansvar , och område C , slutligen , som gäller samarbetet mellan olika regioner i medlemsstaterna eller tredje land , med hjälp av erfarenheter från område A och B , samt samarbete inom forskning och teknisk utveckling , ett ämne som skall fastställas tillsammans med Europeiska kommissionen , som ansvarar för genomförandet .
Det nya Interreg-programmet beaktar man i den form det överlämnats till oss de behov som uppstår genom utvidgningen till länderna i Central- och Östeuropa och till öregionerna och de yttersta randområdena .
Kommissionen föreslår att vi skall fördela Interregs resurser enligt följande : mellan 50 och 80 procent till område A , 6 procent till område C och skillnaden , dvs. mellan 14 och 44 procent , till område B. Europeiska kommissionen fastställer förteckningen över stödberättigade regioner inom område A och B och stöder sig huvudsakligen på kartan över stödberättigade regioner under föregående programplaneringsperiod .
De yttersta randområdena kan åtnjuta stöd inom område B. Kommissionen upprättar en ofullständig förteckning över prioriterade områden och stödberättigade åtgärder för område A , men en fullständig förteckning när det gäller område B. Kommissionen förbehåller sig rätten att senare föreslå frågor som den anser viktiga för utbyte av erfarenheter och förstärkt samarbete mellan regioner inom område C. Förfarandet för att anta programmen fastställs genom den allmänna förordningen om strukturfonderna .
Förslagen upprättas av medlemsstaterna och överlämnas för godkännande till kommissionen , som kontrollerar att de överensstämmer med de allmänna riktlinjer som fastställts .
Dessa förslag måste innehålla ett antal beståndsdelar , en överblick över gränsöverskridande eller transnationella strategier och prioriteringar , en beskrivning över de åtgärder som krävs för att de skall kunna genomföras och en vägledande finansieringsplan .
Jag hör till den stora majoritet av parlamentsledamöter som röstat för att programmet för gemenskapsinitiativet Interreg skall bibehållas .
Jag beklagar att parlamentet inte informerats om utvärderingen av det tidigare programmet - vilket skulle ha gjort det möjligt att göra de nya åtgärderna optimalt effektiva , men jag vet hur svår denna åtgärd är - jag beklagar också att tidsplanen varit extremt kort , eftersom texten granskades i utskottet den 24 november och 26 januari , och jag beklagar också att vare sig de representativa regionerna eller regionala organisationerna fått möjlighet att delta i utarbetandet av programmet .
Genom att främja ett gränsöverskridande samarbete mellan länder eller regioner är detta tvärgående instrument själva inkarnationen av en europeisk regionalpolitik som främjar en harmonisk och balanserad politik för fysisk planering inom gemenskapen .
Fru talman , ledamöter , kommissionärer !
Vid konferensen om landsbygdens utveckling i Cork 7-9 november 1996 klassificerades landsbygdsutveckling som en av Europeiska unionens prioriterade frågor eftersom den är väsentlig för jordbruket , för att uppehålla och kontinuerligt utveckla det , för att ge jordbrukarna nödvändig infrastruktur och service , för en större respekt för miljön och en högre livskvalitet , för diversifiering och skapandet av arbetstillfällen .
Därför anser vi att det fordras en integrerad utvecklingspolitik för alla unionens landsbygdsområden , med följande delområden : ett integrerat och sektorsövergripande synsätt , en förenkling av de administrativa rutinerna , ett utvidgat partnerskap mellan de europeiska institutionerna och nationella och lokala aktörer och ett skydd för miljön .
I programdokumentet Agenda 2000 från 1998 anger kommissionen två huvudprinciper som grund för politiken för landsbygdsutveckling : erkännandet av att jordbruket har många funktioner och behovet av en integrerad strategi för de landsbygdsområden som är under utveckling .
Med denna första princip vill man skapa ett nytt förbund mellan jordbrukaren och samhället genom att göra jordbrukaren till landsbygdens vårdare och tillse att samhället är berett att stå för den miljöservice som fordras för att värna om landsbygdens rekreationsvärde .
Den andra principen grundar sig på konstaterandet att numera en stor del av arbetstillfällena på landsbygden finns utanför den traditionella jordbrukssektorn .
Därför måste man införa ett heltäckande utvecklingsprogram i vilket politiken för landsbygdens utveckling integreras med den sektoriella jordbrukspolitiken : landsbygdsutvecklingen blir därigenom en pelare inom gemenskapens jordbrukspolitik .
Gemenskapens initiativ Leader lanserades 1991 för att främja en ny syn på landsbygdens utveckling , nedifrån och upp , och för att diversifiera åtgärderna genom att de anpassas till de lokala behoven .
Målsättningarna var : att förbättra landsbygdsområdenas utvecklingspotential genom att luta sig mot lokala initiativ , att verka för kunskapsinhämtning inom området landsbygdsutveckling och att sprida denna kunskap till andra landsbygdsområden .
Leader I var inriktat på de landsbygdsområden som omfattades av strukturfondernas mål 1 och 5b .
217 lokala aktionsgrupper deltog i programmet som hade en budget på 1 155 miljoner euro .
Leader II-programmet från 1994 till 1999 - som vi tyvärr ännu inte har en total utvärdering av - hade större omfattning än Leader I. Bidragsmottagarna bör ha varit fler än 800 enheter och avsatta medel efter resursfördelning bör ha överstigit 4 000 miljoner euro .
I oktober 1999 beslöt Europeiska kommissionen mot bakgrund av framgångarna med Leader I och II att förlänga detta initiativ .
För perioden 2000-2006 är tyvärr bara totalt 2 020 miljoner euro avsatta , och en ungefärlig uppdelning mellan medlemsstaterna har gjorts .
Initiativet Leader + skiljer sig från de föregående faserna eftersom denna gång alla landsbygdsområden kan få del av medlen .
Dessutom är det mer ambitiöst och avpassat till de utmaningar landsbygden måste klara .
De viktigaste förändringarna gäller följande aspekter : alla landsbygdsområden kommer att kunna utnyttja Leader + , kriterierna för att välja ut lokala åtgärder blir strängare , de lokala utvecklingsplanerna kommer att läggas in som prioriterade frågor och integreras med hjälp av informationsteknologi , förbättring av livskvalitet och uppvärdering av lokala produkter .
Jag uttrycker alltså min uppskattning av att initiativet fortsätter eftersom det , som jag sade , betonar innovativa utvecklingsstrategier och eftersom det är mer ambitiöst , även om behovet kvarstår att göra kriterierna för vilka områden som omfattas mer flexibla så att man inte straffar varken landsbygdsområden med hög koncentration eller landsbygdsområden med låg koncentration .
Jag anser att nätverkssystemet för utbyte av information och kunskap och för genomförande av gemensamma projekt för olika områden inom unionen är avgörande , och jag påminner om att om det skall kunna förverkligas fullt ut måste man bland annat dra nytta av alla redan befintliga instrument , såsom carrefour .
Jag instämmer i kommissionens åsikt att en lösning av det totala stödet är att föredra , men jag insisterar dock på att redovisningskraven på de nationella och regionala förvaltningarna måste fastställas exakt och ingående .
Jag beklagar att Leader , liksom de tre andra initiativen , framläggs för parlamentet så försenat och den försening detta i sin tur medför för hela förfarandet .
Slutligen bekymrar det mig att det avsatta beloppet är så litet , om man dessutom tar med i beräkningen att programmet denna gång är öppet för alla unionens områden och kommer att gälla ett år längre än föregångaren Leader II .
Jag tackar kommissionens tjänstemän för deras tillmötesgående och samarbetsvilja och kollegerna i utskottet för jordbruk och landsbygdens utveckling för deras bidrag i form av ändringsförslag . .
( DE ) Fru talman , ärade kolleger !
Mitt Equal-betänkande har karaktären av ett yttrande inom ramen för rådfrågningsprocessen för ett nytt gemenskapsinitiativ , vars mål det är att få till stånd ett transnationellt samarbete för att främja nya metoder för bekämpandet av diskriminering och ojämlikheter av alla slag på arbetsmarknaden .
Betänkandet blev mycket kostsamt eftersom det även inbegriper yttranden från fyra andra utskott - från utskottet för industrifrågor , utrikeshandel , forskning och energi , utskottet för regionalpolitik , transport och turism , utskottet för kvinnors rättigheter och jämställdhetsfrågor samt utskottet för rättsliga frågor och den inre marknaden .
Detta gemenskapsinitiativ är en efterföljare till de två föregångarna Adapt och Employment och förfogar över en betydligt mindre budget , nämligen runt 2,8 miljarder euro .
Initiativet slår in på en helt ny väg , nämligen för att ta fram innovativa sysselsättningsmodeller för transnationella utvecklingspartnerskap på geografisk eller sektoriell nivå .
Avsikten är tydlig : det skall utvecklas riktade projekt på transnationell nivå , projekt som orienterar sig efter de sysselsättningspolitiska riktlinjerna , dvs. sysselsättningsförmåga , företagaranda , anpassningsförmåga samt lika möjligheter för alla .
Denna målsättning skall verkligen välkomnas , och den finner gehör även i kammaren .
Equal skall härutöver mynna ut i de nationella sysselsättningsprogrammen samt genom dessa åtgärdsprogram möjliggöra kontroll av införlivandet .
Detta är ett viktigt gemenskapsinitiativ , som tillsammans med de tre andra initiativen Urban , Leader och Interreg finansieras genom strukturfonderna .
Jag har i rapporten försökt reducera de våldsamma förvaltningskostnaderna samt utforma starten på partnerskapet för utveckling något mer öppet och flexibelt .
Jag anser att det tekniska stödet är nödvändigt , men på grund av problemen med de tidigare byråerna för utbyte av information om tekniskt bistånd skall det inte bli något nybildande av dessa byråer innan parlamentets resolution föreligger , och därmed skall förhindras att det politiska ansvaret läggs över på tekniskt bistånd .
Men icke desto mindre är det tekniska biståndet nödvändigt .
Särskild uppmärksamhet skall även riktas mot spridningen av resultaten och mot det ömsesidiga lärandet genom best practice och mainstreaming .
Det har varit min strävan att kunna garantera att betänkandet får ett så brett stöd som möjligt .
Detta har gjort att antalet ändringsförslag har minskats - från över 100 i utskottet till 22 för plenum - och det har sålunda även blivit möjligt att finna talrika kompromisser .
I frågan om asylsökande har det likaledes gjorts en kompromiss .
För att vi även skall kunna utforma detaljerna här ber jag dock , fru talman , att omröstningen om Equal-betänkandet genomförs först på onsdag i stället för i morgon .
Det är viktigt för mig att gemenskapsinitiativet kan köras igång i tid , att betänkandet får ett övertygande stöd så att kommissionen också manas att ta hänsyn till Europaparlamentets konstruktiva förslag , för anslagen till Equal har hållits tillbaka av Europaparlamentet just för att ledamöternas invändningar skall komma till uttryck i detta gemenskapsinitiativ .
Därför är det också befogat att parlamentet insisterar på att ämnesprioriteringarna skall kunna ändras först efter att parlamentet har hörts på nytt .
Equal skall , och det är min bestämda avsikt , göra rättvisa åt sitt namn .
Genom det skall alla eftersatta grupper i Europeiska unionen erbjuda samma chanser .
Det skall förhindra att samhället faller isär .
Det skall hindra utslagningen från att vara en del av vardagen .
Alla skall erbjudas möjligheten att dra fördel av ett gemensamt initiativ , oavsett hur gamla eller av vilket kön de är och varifrån de kommer .
Detta är min avsikt , och jag ber om ett övertygande stöd för betänkandet i kammaren !
Fru talman !
Det är i sig självt en prestation att vi har denna debatt om gemenskapens nya stadsmiljöinitiativ inom Urban-programmet , och det är en prestation att jag är här i kväll , eftersom Air France ställde in mitt flyg som skulle gå kl .
14.10 - men jag är här !
För bara ett år sedan när kommissionen utarbetade sina förslag kring Agenda 2000 skar man ned stadsmiljöinitiativet .
Ändå visste vi i egenskap av politiker att det fanns en underström av stöd för en fortsättning av detta initiativ under år 2000 .
Parlamentet kan därför ta åt sig äran för att ha genomfört en framgångsrik påtryckningskampanj för att få tillbaka Urban-programmet på dagordningen och få kommissionen och rådet att göra en kovändning .
Stadsmiljöpolitiken har alltid varit högt prioriterad inom EU : s politik .
I min medlemsstat , t.ex. , håller vi på att utveckla ett strategiskt förhållningssätt genom en vitbok och en statlig stadsmiljögrupp håller på att undersöka de problem som finns i stadsmiljön .
I ett läge där 80 procent av befolkningen i Europa bor i stadsområden , är det rätt och riktigt att vi hjälper våra mest eftersatta samhällen att ta itu med de alltför bekanta problemen med förfall , social utslagning , arbetslöshet , kriminalitet , drogberoende och alla de problem som har samband med detta .
I min hemregion , t.ex. , i Manchester , har stadsmiljöinitiativet inom Urban-programmet blivit en enorm framgång .
Medel från programmet har investerats i ett av de mest förfallna stadsområdena i Förenade kungariket , Moss Side .
" The Millennium Youth Park " projektet hjälper till med att få unga personer intresserade av att rusta upp sitt eget grannskap och förutom stöd till mindre företag och socialpolitik , börjar vi se en återhämtning inom detta mycket eftersatta stadsområde .
Arbetet med denna Urban-dagordning togs sedan till andra delar av samhället med en aktiv kommunikations- och offentlighetskampanj på lokala stormarknader och berömda brittiska pubar .
Det är denna typ av bra åtgärder som vi också vill skall utvidgas till hela EU när det rör kommunikation och offentlighet .
Vad gäller de särskilda riktlinjer som styr initiativet , är de flexibelt definierade för att ge utrymme för lokal och regional mångfald .
Vi håller med om att de bör vara vägledande till sin natur och låta en maximal flexibilitet se till att vi uppnår specifika programmål .
I utskottet förespråkar vi inte en minskning av antalet till 50 .
Vi förespråkar en allmän minskning , men vi anser inte att den godtyckliga siffran 50 är den viktigaste faktorn .
Vi borde i stället satsa på högkvalitativa projekt som kan fungera som en katalysator för förändring och förnyelse , som kan dra till sig investeringar rörande lån och riskkapital och åstadkomma en multiplikatoreffekt .
Medlemsstaterna bör därför kunna föreslå ett skäligt antal områden inom det finansiella taket för sina anslag .
Vid angivandet av lokala Urban-program , måste vi verkligen ta hänsyn till lokala indikatorer och lokal statistik om eftersatthet och hälsotillstånd för att vi skall kunna ta itu med de värst drabbade områdena på ett mer effektivt sätt .
I Förenade kungariket är det lokala eftersatthetskriteriet ett mycket bra exempel på en allmänt använd standard och statistik till hjälp för att bestämma inte bara stödprogram inom EU , utan också nationella och regionala stödprogram .
Detta måste börja användas som ett instrument och en resurs , som ett komplement till EU-kriterierna .
Jag vill be er att ta hänsyn till lokala indikatorer för att hjälpa oss med detta .
Våra mest eftersatta stadsområden står inför en överväldigande mängd problem : Hög arbetslöshet och ofta mycket dåligt betalda och osäkra jobb , fattigdom och social utslagning .
Dessa problem förvärras ofta genom dåligt hälsotillstånd , dåliga bostäder och en kultur där drogberoende ingår .
Det är därför vi har fått instabila samhällen som genomsyras av kriminalitet , narkotikahandel och gäng .
Detta är alltför välbekant i många av våra stadsområden .
Alla dessa komplexa problem undergräver livskvaliteten för de stadsboende , fast möjligheten finns i dessa områden att skapa tillväxt och välstånd .
Detta är återigen skälet till varför jag i mitt betänkande har poängterat att åtgärder i samband med Urban-programmet inte bara bör tillhandahålla en helhetslösning till ett enda problem : Dessa områden lider inte av enstaka problem .
Samhällena i stadsområdena bör i stället uppmuntras till att lägga fram integrerade handlingsplaner som kan hjälpa till med att lösa deras specifika stadsrelaterade problem , genom att använda EU-resurser som ett komplement till lokala åtgärder .
Jag skulle vilja se att dessa åtgärder utökades till att omfatta hälsofrågor och åtgärder mot diskriminering , som fastställts i Amsterdamfördraget .
Gemenskapsinitiativet innebär gemenskapsengagemang .
Några av de mest aktiva och engagerade krafterna för förändring inom våra stadsområden är de personer som bor där .
Vi måste uppmuntra dem att delta i utformningen och slutförandet av projekt inom dessa program .
Den tidtabell som föreslagits av kommissionen är därför mycket ambitiös .
Det är bättre att ha kvalitetsprojekt med ett aktivt deltagande av gemenskapsgrupper , än att ha projekt som slutförs enligt tidtabell men utan lokalt deltagande .
Kommissionen måste naturligtvis se till att det råder fullständig öppenhet rörande de urvalskriterier som används för de nya programinitiativen , men den måste också redovisa vilka rådgivningsnätverk som används för utbytet av bästa metoder .
Detta är viktigt när det rör öppenhet och nätverkens övergripande effektivitet .
Låt mig till sist betona att vi behöver lokalt engagemang för att kunna ta itu med de problem som det postindustriella samhället står inför .
Vi måste använda oss av de arbetslösas inneboende kraft , ungdomarnas för litet använda färdigheter och de äldres erfarenheter för att kunna lösa dessa problem .
Vi skall då kunna ersätta fattigdom , beroende och främlingsskap med rättvisa , initiativkraft och deltagande .
Detta kommer att hjälpa oss att återställa EU : s trovärdighet och medborgarnas tro på att Europeiska unionen kan få till stånd lokala åtgärder för att lösa lokala problem . .
( IT ) Herr talman !
Som föredragande McCarthy redan har påmint om kan Urban verkligen betraktas som en seger för Europaparlamentet som en följd av den debatt som pågick förra året om reformering av förordningarna .
Som har sagts är syftet med Urban att främja innovativa strategier till förmån för en ekonomisk och social nylansering av stadsområdena , också mot bakgrund av att 80 procent av Europas befolkning är koncentrerad till städerna .
Att skapa en positiv stadsmiljö ur socialpolitisk synvinkel innebär att förverkliga en politik som syftar till att skapa varaktiga arbetstillfällen , att bekämpa fattigdomen , att vidta åtgärder till förmån för låginkomsttagare , äldre och barn , etnisk och rasmässig integration , bättre möjligheter till delaktighet , en profilerad hälso- och sjukvårdspolitik som omfattar åtgärder för att förebygga drogberoende liksom en samordnad brottsförebyggande politik .
Kommissionen tar i sitt meddelande hänsyn till behovet av angreppssätt som omfattar ett helt spektrum av ekonomiska och sociala infrastrukturåtgärder .
Emellertid måste man komma ihåg att det förutom Urban finns flera andra gemenskapsinstrument på det sociala området : innovativa åtgärder enligt Europeiska socialfondens artikel 6 , pilotprojekt - framför allt den nya förberedande satsning på " Lokala sysselsättningsinitiativ " , som Europaparlamentet nyss införde i och med budgeten för 2000 - initiativen Equal och Interreg liksom mainstreaming av socialfonden .
Som utskottet för sysselsättning och socialfrågor understryker i sitt yttrande måste alltså kommissionen ta hänsyn till synergieffekter i detta sammanhang och samtidigt undvika dubbleringar inom de finansierade projekten .
Samtidigt som vi å ena sidan anser det nödvändigt att styrkommittéerna säkerställer att de olika insatserna är inbördes konsekventa och kompletterar varandra , uppmanar vi å den andra sidan kommissionen att öka informationsutbytet och samordningen mellan de avdelningar som berörs .
En sådan samordning är inte det enda som är viktigt , utan även utbytet och spridandet av erfarenheter och god praxis måste vara viktigt , vilket vi påpekar i vårt yttrande .
Herr talman !
Betydelsen av detta initiativ blir allt större allt eftersom de ekonomiska och sociala problemen förvärras i Europas städer och allt eftersom invånarna i städerna känner sig allt med fjärmade från sina städers eller förorters förvaltning .
Till denna situation kommer de sociala omstruktureringarna till följd av utvidgningen av Europeiska unionen att komma till , och följaktligen måste vi i god tid ombesörja våra städers ekonomiska förnyelse och sociala sammanhållning .
Dessa problem måste för övrigt bemötas även med tanke på städernas stora inflytande på de kringliggande regionerna , liksom även med tanke på deras historiska och kulturella roll .
För att våra ansträngningar skall lyckas , krävs det emellertid att alla medborgare engagerar sig och deltar samt att de mindre aktiva samhällsgrupperna och de grupper som drabbas särskilt hårt av den ekonomiska och sociala krisen aktiveras .
Och här vill vi betona nödvändigheten av att kvinnorna , eller de aktörer som företräder kvinnorna , på ett balanserat sätt deltar i planeringen och genomförandet av Urban-initiativets program .
Vi i utskottet för kvinnors rättigheter och jämställdhetsfrågor betonar även nödvändigheten av att finansiera infrastrukturer som gör det lättare för kvinnorna att vara yrkesverksamma , huvudsakligen med avseende på en harmonisering av yrkes- och familjeansvaret , och bredare infrastrukturer som främjar generationernas solidaritet , den sociala solidariteten .
Om detta initiativ genomfördes på ett effektivt sätt , skulle det kunna få en multiplikatoreffekt , eftersom det skulle kunna stimulera till liknande åtgärder på regional och lokal nivå .
Initiativets politiska betydelse skulle då bli ännu större , eftersom kvinnorna behöver känna påtagliga resultat av den europeiska politiken i sina vardagliga liv. ån utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor .
( DE ) Herr talman !
Vi har i vårt utskott välkomnat det faktum att kommissionen har föreslagit att Urban-programmet skall prioritera en bättre integrering av lokala gemenskaper och etniska minoriteter liksom höjningen av säkerheten och förebyggande åtgärder mot kriminalitet .
Vi har i utskottet ansett det nödvändigt att ett ekonomiskt och socialt återupplivande av stadsområden åtföljs av en atmosfär med tolerans gentemot minoriteter , så att åtgärder avsedda att minska rasism och främlingsfientlighet blir ett integrerat inslag i de program som skall finansieras inom ramen för Urban .
Vi har ansett att en central uppgift när det gäller återupplivandet av stadsområden är att höja medborgarnas känsla av trygghet och därmed att bekämpa vardagskriminaliteten i städerna .
Utskottet har konstaterat att en nytänkande och effektiv kriminalitetsbekämpning liksom förebyggandet av kriminalitet kräver åtgärder som differentieras på kommunal nivå - hit hör att förebyggandet av kriminalitet tas med i stadsplaneringen , åtgärder för att förebygga ungdomsbrottslighet , återanpassning av förbrytare liksom modeller för ett verkningsfullt samarbete mellan olika aktörer på lokal nivå , t.ex. polis , rättsväsende eller sociala instanser .
I utskottet har vi enhälligt ställt oss bakom rekommendationen , eftersom vi var mycket angelägna om att just Urban - som i tidigare skeden har varit ett så framgångsrikt gemenskapsinitiativ - får en fortsättning , för vi utgår ifrån att vi endast med hjälp av dylika program inom Europeiska unionen kommer att lyckas förverkliga en fredlig samexistens på sikt för alla invånare i Europeiska unionen .
Det är av den anledningen som vi varmt välkomnar denna typ av program. ättning och socialfrågor .
( DE ) För det mest omfattande av de fyra gemenskapsinitiativen , nämligen Interreg III , vill jag föra fram önskemålen från utskottet för sysselsättning och socialfrågor .
Det måste finnas möjlighet att satsa stort även på sociala åtgärder när det gäller Interreg III .
Med tanke på att 50 procent av arbetslösheten i unionen till väsentliga delar är strukturellt betingad och med tanke på den särskilt känsliga situationen i gränsområdena - jag pekar endast på möjliga oönskade migrationsrörelser - är detta inte bara förnuftigt , utan nödvändigt .
Nu tycks också de stödåtgärder som anförs i bilaga II till programinriktning A vara lovande i detta hänseende .
Men i kommissionens meddelande saknas det faktiskt helt och hållet bestämmelser för medlemsstaterna som omfattar dessa integrerade satsningar på social- och sysselsättningspolitiska aspekter .
Därför vill jag särskilt betona ett ökat insättande av yrkesutbildningsåtgärder , i synnerhet i områden med hög långtids- och ungdomsarbetslöshet .
Inriktning B bör likaledes vara öppen för sysselsättningspolitiska stödåtgärder , speciellt i samband med strategin för att föra fram medlemskandidaterna .
När det gäller de sysselsättningspolitiska åtgärderna ser jag det rent generellt som en nödvändighet att den gemensamma samarbetskommittén tillsätts regionalt därför att närheten och den nödvändiga sakkunskapen som rör dessa åtgärder bara finns på regional nivå och därför att det skall förhindras att åtgärderna blir verkningslösa .
Att förvaltningskostnaderna för Interreg III - som jag ser det - fortfarande är för höga kan vi alltid kritisera , det måste vi också hela tiden göra , även om jag nästan börjar tro att detta är oundvikligt i kommissionens stödprogram .
Jag vill dock påpeka att det är ödesdigert just här .
Just vad gäller sysselsättningspolitiken bör vi eftersträva så enkla åtgärder som möjligt för att den sociala dimensionen i Europeiska unionen återigen skall ges den tyngd som den förtjänar .
Herr talman !
Utskottet för regionalpolitik , transport och turism tittade bl.a. på meddelandet om Leader + och beslutade att stödja decentraliseringsprocessen i hanteringen av åtgärder .
Man ansåg att en sådan process kan vara effektiv om man uppfyller två villkor : att de lokala aktionsgrupperna är representativa för lokalsamhällets allmänna intressen och att kommissionens kontrollmekanismer används för att undvika att de territoriella och lokala myndigheterna använder medel från Leader + för att bibehålla organisationer och civila grupper vinklade till myndigheten .
Det begärs att man i de organ som fattar beslut om projekten garanterar en likvärdig representation av tre komponenter : de politiskt valda och offentliga myndigheter , företagen och de ekonomiska parterna , samt arbetsmarknadens parter , inklusive fackföreningar och frivilligorganisationer .
Särskilt understryks att det skall vara en jämn könsfördelning i alla dessa organ .
Man understryker dessutom att huvudsyftet är att främja strategier för en hållbar utveckling , vars positiva effekter skulle sträcka sig över ett bredare geografiskt område än själva lokalsamhället , och man anser det således vara lämpligt att projekten innefattas i utvecklingsprogrammen , inklusive mål 1 och 2 samt i planerna för den fysiska planeringen i de regioner och länder där de lokaliseras .
Man gläds åt att Leader + kan användas i alla landsbygdsområden i unionen , men man beaktar dock att det är nödvändigt med en koncentration av gemenskapsresurserna till de mest missgynnade regionerna för att underlätta den socioekonomiska sammanhållningsprocessen i unionen , utan att de statliga myndigheterna styr dessa medel mot syften som inte har med sammanhållningen att göra .
Utskottet är av den uppfattningen att man för de projekt som finansieras inom ramen för åtgärd 1 borde värdera potentialen för en endogen utveckling , som i synnerhet stöds på lokala traditioner , tekniker och vanor , på specifika produktioner och på en hållbar energiutvinning .
Utskottet stöder kommissionens förslag att koncentrera åtgärderna till ett reducerat antal valda områden och är av den uppfattningen att med hänsyn tagen till de olikheter som finns i många samhällen på landsbygden skall det demografiska minimitaket för att välja ett projekt minskas till 10.000 invånare .
Man anser att det är nödvändigt att samordna utvecklingsmålen och mekanismerna för hantering av åtgärderna 2 och 3 som finansieras av Leader med övriga åtgärder som finansieras med hjälp av andra gemenskapsprogram för samarbete och interregionala och internationella partnerskap , som Interreg , Sapar , Phare , Tacis och Meda inom samma områden . .
( IT ) Herr talman !
Jag skall tala om Equal-betänkandet i två minuter för utskottet för kvinnors rättigheter och jämställdhetsfrågor och sedan i två minuter för socialistgruppen i utskottet för sysselsättning och socialfrågor .
Gemenskapsinitiativet Equal , vars mål är att verka för nya instrument som skall bekämpa alla former av diskriminering och ojämlikhet , behandlades mycket ingående i utskottet för kvinnors rättigheter och jämställdhetsfrågor ur aspekten kvinnodiskriminering .
Detta beror på att könsbaserad diskriminering är strukturell och horisontell och att utskottet för kvinnors rättigheter och jämställdhetsfrågor - mot bakgrund av att kvinnorna inte utgör en minoritet utan mer än hälften av världens befolkning - anser att det kanske var fel att ta med könsbaserad diskriminering bland all annan diskriminering .
Vi anser att det hade varit bättre att lägga in den könsbaserade diskrimineringen i ett särskilt kapitel i fördraget om lika möjligheter för män och kvinnor , som en logisk konsekvens av den nya centrala roll jämställdhet mellan män och kvinnor har fått i fördraget .
När detta är sagt gläder vi oss ändå åt kommissionens förslag och hävdar att jämställdhet mellan män och kvinnor bör främjas som en integrerad del i alla de fyra pelarna i sysselsättningsstrategin liksom i sakfrågorna och samtidigt vara en egen särskild pelare .
Vad Equal-föreslagen beträffar anser vi att man i programmen i gemenskapsinitiativen bör göra klar åtskillnad mellan prioriterade åtgärder i syfte att bekämpa könsdiskriminering och andra former av diskriminering och att man bör tillämpa ett angreppssätt som syftar till att införa jämställdhet mellan könen i all gemenskapspolitik , och alltså betonar nödvändigheten av att även verkställa projekt som syftar till att bekämpa inte bara könsdiskriminering utan också att underlätta för människor att förena familje- och yrkesliv .
Mer generellt hade utskottet för sysselsättning och socialfrågor en mycket omfattande debatt om Stenzels betänkande eftersom det angreppssätt han föreslog skilde sig mycket från min grupps .
Vi har bedömt kommissionens förslag som någonting mycket positivt , men ändå försökt finna lösningar som vi kan vara överens om , så att betänkandet kan röstas igenom av en bred majoritet .
Målet var ju nämligen att Europaparlamentet skulle avge ett yttrande som sedan skulle väga tungt under kommissionens och rådets överväganden .
Vissa punkter var mer känsliga än andra : till exempel partnerskapen , där jag tror att man måste finna en kompromiss för att stärka och stödja kommissionens förslag .
Samtidigt måste man dock be kommissionen om en viss flexibilitet så att man senare kan lägga in andra frågor .
Likaså måste den tekniska servicen och förenklingen finnas med bland de grundläggande punkterna .
Den mest känsliga frågan ur politisk synpunkt var den om de asylsökande .
Jag vill uppehålla mig vid detta ämne några sekunder eftersom vi anser att kommissionens förslag är komplett och positivt .
Vi har lagt ned mycket tid på att hitta en definition av asylsökande eftersom detta är svårt juridiskt sett , men jag tror att vi nu har uppnått en kompromiss med föredraganden - åtminstone hoppas jag det - och att det betänkande parlamentet kommer att rösta om tiger om asylsökande skall ses som ett stöd för kommissionens ståndpunkt från parlamentets sida .
Vi skulle aldrig ha accepterat att parlamentet tog ett steg tillbaka - detta är vår inställning - jämfört med kommissionens förslag , och detta vill jag understryka .
Jag instämmer med föredraganden om att vi bör rösta på onsdag , som hon föreslog , så att vi har tid att hitta alla upptänkliga lösningar för att göra parlamentets betänkande kanske till och med mer avancerat , inte mindre , än kommissionens förslag . .
( DE ) Ärade herr talman , ärade fru föredragande , ärade kolleger !
Innan jag närmare går in på Equal-betänkandet vill jag säga något principiellt om de riktlinjer för sysselsättning som ligger till grund för betänkandet .
De grundläggande målen med en gemensam sysselsättningspolitik för EU har där fastställts till att gälla bland annat sysselsättningsförmåga , företagaranda och anpassningsförmåga .
Dessa mål syftar uppenbarligen till att göra arbetstagarna så nyttiga och exploaterbara som möjligt för näringslivet .
Ett försök att verkligen avveckla diskriminering på ett effektivt och långsiktigt sätt skulle emellertid behöva ha människors självbestämmande som mål .
Först då handlar det inte längre endast om ekonomisk användbarhet , utan om ett jämlikt sätt för människor att gestalta sina liv .
Likväl har Stenzels betänkande utvecklats bra , åtminstone det som rör de fastställda riktlinjerna .
Alla asylsökande och flyktingar skall uttryckligen omfattas av programmet , vilket emellertid borde vara en självklarhet .
Ändå har de konservativa i utskottet röstat emot detta .
Till dessa personer har jag en fråga : Är målet med er politik att marginalisera människor ?
Vad är det för idé som ligger bakom att förvägra människor arbete när de vill arbeta ?
Står inte det i rak motsats till riktlinjen " sysselsättningsförmåga " ?
Det är också värt att nämna att det här handlar om ett mainstreaming-program , för betänkandet är förenat med vissa brister .
Sålunda betonas särskilt aspekten att kvinnor skall beredas bättre möjligheter på arbetsmarknaden genom att fler förskolor skall byggas .
Den som låter männen klättra ostört uppför karriärstegen och enbart bekymrar sig om daghemsplatser utan att bekämpa den ojämna fördelningen av det reproduktiva arbetet , han och dessvärre även hon har inte förstått vad mainstraming är !
Herr talman , ärade damer och herrar !
Utskottet för regionalpolitik , transport och turism har vid de avslutande överläggningarna enhälligt , dock med en nedlagd röst , godkänt föreliggande yttrande om Equal-betänkandet .
Detta placerar jag medvetet först i min redogörelse för att tydliggöra att det faktiskt föreligger en motsättning mot det ansvariga utskottet för sysselsättning .
Att samtliga grupper har godkänt yttrandet kan förklaras av de slutsatser som är ägnade att koppla samman regional- och transportpolitiska frågor liksom turismfrågor med bekämpningen av diskriminering och ojämlikheter av alla slag på arbetsmarknaden .
Ledamöterna i utskottet för regional ser naturligtvis även en rad kritiska moment i kommissionens förslag , för det första har exempelvis den tematiska orienteringen för utvecklingspartnerskapens agerande inte fastställts i tillräcklig utsträckning ; för det andra återstår det fortfarande för kommissionen att utarbeta strikta urvalskriterier för utvärderingen av projektförslagen ; för det tredje befarar man för höga förvaltningstekniska kostnader för projektledningen via kommissionen liksom instanserna för det tekniska biståndet .
Därför skall en övre gräns dras för förvaltningsuppgifterna .
Utskottet har dragit slutsatser av dessa kritiska anmärkningar .
Särskild vikt lägger vi vid kopplingen mellan skapandet av nya arbetstillfällen för socialt missgynnade och utslagna personer , inom turismen såväl som inom de små och medelstora företagen , och stödet för bildandet av små och medelstora företag med hänsyn till den nödvändiga ekonomiska strukturförändringen .
Sammanflätningen av aktiviteterna inom gemenskapsinitiativen och de europeiska sysselsättningsinitiativen är ett grundläggande krav och en avgörande förutsättning för att Equal-programmets olika uppgifter skall kunna fullgöras .
Vi stöder eftertryckligen det innovativa försöket att bilda internationella utvecklingspartnerskap och att organisera utbytet av erfarenheter på europeisk nivå som en integrerad beståndsdel i Equal-programmet .
Den speciella målsättningen att nå europeisk framgång lyfter upp det regionala samarbetet till europeisk nivå samtidigt som samarbetet mellan de mest skilda regionala aktörer bibehålls .
Detta är bra , och därför har vi också rekommenderat det .
Herr talman , mina damer och herrar , kära kolleger !
Det har redan påpekats i dag att det första Urban-initiativet var entydigt framgångsrikt .
Att detta initiativ nu skall få en fortsättning som Urban II , om än med minskade anslag , har vi enskilda engagerade ledamöter av parlamentet att tacka för , särskilt - så vitt jag som ny ledamot av parlamentet förstår - föredraganden fru McCarthy som jag därför vill tacka så hjärtligt för hennes insats och naturligtvis även för hennes betänkande om Urban II .
( Applåder ) Nytt i Urban II-initiativet är att det har inriktats på små städer och stadsdelar .
Detta är viktigt eftersom just små städer ofta har sämre möjligheter att få stödanslag .
Å andra sidan kan det hända att de problem som leder till stort behov av förnyelse gärna koncentreras till just sådana städer och i motsvarande mån får starkt negativa följder .
För att öka de enskilda åtgärdernas effektivitet har antalet projekt för Urban II begränsats till 50 .
Jag tycker det är viktigt att inte hålla stelt på denna godtyckligt satta siffermässiga begränsning utan att överlåta åt medlemsstaterna att avgöra på hur många projekt var och en vill fördela de stödanslag man är berättigad till .
Men det gäller att ge akt på att det just i de små medlemsstaterna ändå inte bara blir stadsdelar i storstäder som kommer i åtnjutande av stödet .
Där vore Urban II bara en droppe i havet , av tvivelaktigt resultat , och det skulle falla platt till marken .
Lika viktigt är det enligt min mening att urvalskriterierna för Urban II inte utvidgas överdrivet , så att de därigenom urvattnas .
Just en strängt avgränsad kriteriekatalog är en förutsättning för att de stödda projekten skall få modellkaraktär och i framtiden kunna överföras på andra problemstäder .
Min egen kommunalpolitiska erfarenhet från en gammal industrialiserad region med många problem gör att jag avslutningsvis vill be er , kära kolleger , om särskilt stöd för två punkter i rapporten , vilka jag vid sidan av de socialpolitiska aspekterna anser vara väsentliga .
För det första : miljöskyddsaspekten är absolut nödvändig för en hållbar stadsutveckling och bör därför vara en generell förutsättning för projektstödet .
För det andra : Förebyggandet och bekämpningen av vardagskriminaliteten i städerna liksom av kriminaliteten kring anskaffandet av droger måste börja på lokal nivå .
Detta är absolut nödvändigt för en ökad urban livskvalitet och måste därför spela en central roll i Urban II-initiativet .
Herr talman , bästa föredragande , bästa åhörare !
Jag tackar föredragandena som på kort tid åstadkommit sakkunniga betänkanden .
I min grupp har man dock kritiserat tidpunkten för utskottets förberedelsearbete .
Betänkandena är försenade , dessutom drevs behandlingen åtminstone i utskottet för regionalpolitik , transport och turism med en stor brådska .
På så vis missade man ett bra tillfälle att debattera resultatet av tidigare program , god praxis och även brister .
Vår grupp betonar i samband med Interreg-programmet den gränsöverskridande verksamheten och i synnerhet det samarbete som sträcker sig utanför unionens gränser .
Viktiga regioner är bland annat Balkan och regionerna vid Adriatiska havet , men enligt min mening bör man inte heller glömma samarbetet med Ryssland .
Vår grupp vill på nytt lyfta upp den praktiska kontrollen av fonderna och framhåller bland annat vikten av en bättre samordning mellan Interreg- , Tacis- , Ispa- och Phare-programmen .
I dag saknas denna samordning , och kommissionen har fortfarande inte lagt fram exakta förslag för att förbättra samordningen .
Vi här i parlamentet förväntar oss att kommissionen så snabbt som möjligt skall lämna en noggrannare redogörelse av frågan inför vårt utskott .
När det gäller det praktiska genomförandet är det av avgörande betydelse att få med sig lokala företag , organisationer och andra aktörer .
Erfarenheten har visat att det i samarbetsprojekten behövs bättre planering , noggrannare uppföljning och genomförande som leder till bättre resultat .
Projekten har ofta stannat halvvägs och effektiviteten försvunnit i förvaltningen och byråkratin .
Man måste också kräva av samarbetspartner att de förbinder sig till projekten och uppfyller sin egen del .
Vår grupp lägger på nytt fram några ändringsförslag som avslogs vid utskottsbehandlingen .
Jag tar här upp Urban-betänkandet där föredraganden i motiveringar på ett förtjänstfullt sätt behandlat det minimibelopp på 500 euro per invånare som ingår i kommissionens riktlinjer .
Det fungerar inte som ett mekaniskt mål utan det måste kunna anpassas efter förhållandena i målområdet .
Detta är en så viktig synpunkt att det måste lyftas från motiveringar till slutsatser .
Herr talman , kära kolleger !
Interreg är en av de mest europeiska av alla strukturfonder .
Här skall projekt stödjas inte bara i en region , i ett land , utan i angränsande regioner i två eller flera länder .
Tyvärr gäller detta endast en del av pengarna , nämligen endast för gränserna inom EU .
Men just de regioner som gränsar till tredje land är de som behöver ett fungerande verktyg för ett gränsöverskridande samarbete .
Förordningen ger sken av att det också skulle förhålla sig så .
Men så förhåller det sig inte .
Det förhåller sig nämligen så att kommissionen inte har ändrat förordningen på flera år , trots att parlamentet kräver detta sedan länge .
För regionerna innebär det i praktiken att det den närmaste tiden återigen degraderas till att likna Västtysklands tidigare stödåtgärder till förfallna områden längs gränsen mot Östtyskland .
Parlamentet har sedan 1996 krävt att en gemenskapsfond bildas för samarbetet med tredje land för att lösa problemen .
Ingenting har hänt !
Man drar ytterligare ut på tiden med problemen , på berörda regioners bekostnad .
Parlamentet kräver på nytt en förbättring och ett gränsöverskridande samarbete , och vi förväntar oss att en gemenskapsfond bildas och att förordningen ännu en gång ändras i samarbete med övriga kommissionärer .
Vi vill ha ett medborgarnas Europa och inte ett byråkraternas Europa !
Herr talman !
En tredjedel av Europeiska unionens pengar stoppas in i fonder för allehanda utvecklingsändamål .
Min grupp anser att det är utmärkt om detta leder till att man arbetar bort eftersatta regioner , städer eller befolkningsgrupper eller att hälsan och miljön förbättras .
Det är en fråga om solidaritet och utveckling .
Men att dela ut alltmer pengar är ingen garanti för att de också används på ett allt bättre sätt .
Kommunerna och regionerna där pengarna hamnar har med tiden fått praktisk erfarenhet .
De konstaterar att det är ytterst svårt att använda pengarna till de ändamål där de allra bäst behövs .
Det brukar för det mesta gå bra med allt som faller under ekonomisk tillväxt och infrastruktur , men det är ofta inte helt säkert att sociala ändamål och miljösyften blir godkända .
Eftersom det råder stor osäkerhet om hur reglerna skall tolkas hyr kommuner och regioner nu in dyra byråer .
Dessa sakkunniga får till uppgift att göra en uppskattning av i vilken grad Europeiska kommissionens tjänstemän är beredda att godkänna planerna .
I vissa fall får jag intryck av att det inte handlar om solidaritet eller om att lösa de mest akuta problemen , utan om att upprätthålla befintliga intressen och om propaganda för Europeiska unionens välsignelser .
Det förefaller som om den viktigaste målsättningen på detta område har blivit att snickra ihop och måla propagandaskyltar där det står att ifrågavarande projekt medfinansieras av Europeiska unionen .
Det är för mycket pengar som går till spillo på propaganda och utredningsbyråer , på överläggningar och kontroll , och mycket pengar går tillbaka till det land som de kom ifrån .
Efter den planerade anslutningen av nya medlemsstater med 100 miljoner invånare , där välfärdsnivån ligger på en tredjedel till två tredjedelar av genomsnittet för dagens medlemsstater i Europeiska unionen , kommer detta slöseri att skapa ännu fler nackdelar .
I utskottet för regionalpolitik , transport och turism var gruppen enade vänstern överens med föredraganden av yttrandet om Leader , Nogueira Román .
Med rätta konstaterade denne att det inte ligger något positivt i att sprida alla dessa medel över alla landsbygdsområden .
I valet mellan innovationsprojekt och att koncentrera pengarna till att bekämpa eftersatthet väljer vi det sistnämnda eftersom detta ger det största bidraget till jämlikhet .
Innovation i områden där det redan går bra ger ju redan avkastning och kommer att äga rum även utan europeiska bidrag .
Ytterligare en punkt att uppmärksamma är risken för maktmissbruk och svågerpolitik inom regionala och kommunala förvaltningar .
Tonvikten ligger på lokala grupper där myndigheter , organisationer och vinstinriktade företag samarbetar .
Diskussionen har handlat om den fördelningsnyckel som skall tillämpas i sammanhanget .
Här har bland annat en variant varit på tal som för tankarna till den nederländska " poldermodellen " , det strukturellt organiserade samarbetet mellan stat , fackförbund och företagarorganisationer .
Låt oss inte glömma bort att val till kommunfullmäktige och regionala församlingar hålls för att företräda hela befolkningen .
Egentligen borde det vara så att dessa organ gör en avvägning och då tar hänsyn till fackföreningsrörelsens och miljörörelsens önskemål .
Min grupp motsätter sig inte att fackföreningsrörelsen och miljörörelsen , vars insatser i samhället vi anser vara viktiga , tilldelas en egen tydlig roll .
Det kan förekomma att deras insatser förbigås på grund av lokala förvaltningar som fungerar kortsiktigt eller som inte fungerar tillräckligt demokratiskt .
Men det faktum att vi nu måste vara rädda för maktmissbruk och svågerpolitik antyder att demokratin tyvärr ännu inte fungerar optimalt .
En invändning är att de valda organens begränsade roll medför att företag får mer inflytande .
Så länge ekonomin inte vilar på demokratiska avvägningar av allas behov i stället för vinstintresset för några få är det tveksamt om demokratin fungerar bättre under inflytande från företagare än under inflytande från kommunfullmäktige .
För oss handlar det om " en människa , en röst " i stället för " en aktie , en röst " .
Herr talman !
Det finns ekonomiska gränser inom Europeiska unionen och vid rådande tidpunkt fungerar den inre marknaden med fri rörlighet för varor , personer , tjänster och kapital helt och fullt .
Men om den inre marknaden skall kunna fungera effektivt och om den gemensamma europeiska valutan skall bli framgångsrik , är det viktigt att alla regioner i Europa - det finns över 100 - kan konkurrera ekonomiskt inom denna mycket utmanande miljö .
Vissa områden i Europeiska unionen är ekonomiskt sett mycket starka och överskrider mycket tydligt den genomsnittliga inkomsten per capita .
Det finns fattiga regioner i unionen som måste få stöd från gemenskapen för att förbättra strukturerna hos sina ekonomier , så att de kan konkurrera inom Europeiska unionens struktur .
Om vi tittar på EU : s budgetplan mellan 1989 och 1993 , och 1994 och 1999 , är det därför vi kan konstatera att en så stor andel av EU : s budget avsattes för förvaltningen av Europeiska regionala utvecklingsfonden och Europeiska socialfonden .
Det finns dubbla problem som fortfarande återstår för många europeiska regioner : För det första har vi bristen på lämplig infrastruktur vad gäller vägar , vattenreningsanläggningar och transportnät i detta sammanhang ; för det andra har vi behovet av att få igång initiativ för att bekämpa ungdoms- och långtidsarbetslöshet , som är ett ständigt socialt problem i många stads- och landsbygdsområden i Europa .
Det måste alltid finnas ett engagemang för att se till att vi inte bara bygger ett städernas Europa .
Vi måste se till att det sätts igång sysselsättningsskapande initiativ som främjar sysselsättningen inom sektorn för små och medelstora företag , även på den europeiska landsbygden .
De huvudsakliga aspekterna av debatten denna kväll har samband med funktionen hos gemenskapsinitiativen , dvs. de nya Interreg III- , Equal- och Leader + -initiativen .
Mellan dessa tre program måste det finnas en tydlig demonstration av EU : s engagemang för främjande av en gränsöverskridande utveckling , kampen mot problemen i samband med långtidsarbetslöshet och stöd till program för landsbygdsutveckling .
Herr talman !
Det finns en hel del städer i Europeiska unionen som har att kämpa med det underläge de befinner sig i .
Det finns inte alltid tillräckligt med medel tillgängliga inom medlemsstaterna för att ta itu med detta på ett effektivt sätt .
Därför är det meningsfullt att Europeiska unionen fortsätter att stödja medlemsstaterna och , om så behövs , ger kompletterande stöd inom ramen för Urban .
Kommissionens förslag beträffande Urban innehåller en nedskärning för de kommande sju åren , både i fråga om gemenskapsbudgeten och antalet gynnade områden .
Jag tvingas i likhet med kollega McCarthy konstatera att antalet områden har skurits ned på ett ganska drastiskt sätt .
Det vore önskvärt med en viss frihet för medlemsstaterna att inom en viss budget själva bestämma antalet projekt .
Vad budgeten beträffar så består Urban som sagt av stöd och komplettering till den nationella politiken .
Om så behövs för att generera extra medel är det enligt min uppfattning också helt logiskt att i första hand vända sig till medlemsstaterna och privata finansiärer .
De gröna kan därför inte räkna med vårt stöd för ändringsförslag 2 , vilket de inte heller fick under utskottssammanträdet .
Dessutom anser jag att stöd till en stad eller en trakt , i synnerhet där det handlar om gemenskapsbidrag , måste ha en stimulerande effekt .
Strukturellt stöd skulle leda till bidragsberoende .
På det sättet skjuter vi över målet .
Slutligen bara en allmän kommentar om Interreg .
Stöd till gränsöverskridande projekt skall enligt min uppfattning endast beviljas om regionerna verkligen önskar att få detta .
Vid genomförandet av projekten är det också viktigt att de inte står i strid med den allmänna gemenskapslagstiftningen .
Enligt revisionsrättens rapport för år 1998 är det inte någon inbillad risk .
Det är också anledningen till vårt ändringsförslag för att förebygga motstridigheter mellan allmän politik och konkreta projekt .
Jag tar mig friheten att först av allt uttrycka min bestörtning över de 14 rådsrepresentanternas förhastade fördömande av Österrike .
Herr talman , kära kolleger !
Reformen av strukturfonderna leder till att gemenskapsinitiativen koncentreras till sammanlagt fyra .
Jag välkomnar fortsättningen på och den framskjutna placeringen av Interreg .
Dock orsakar förseningen av direktivförslaget ett par problem .
Regionerna inkluderades inte i tillräcklig utsträckning i förberedelserna till direktivet , trots att det under diskussionen om reformen av strukturformerna ofta krävdes att så skulle ske .
Det saknas en direkt övergång mellan Interreg II och III , vilket i praktiken drar med sig osäkerhet i planeringen och luckor i finansieringen .
Det är synd , för det äventyrar verkligt meningsfulla projekt .
Vid genomförandet av Interreg måste samordningen och synkroniseringen med övriga berörda finansinstrument tryggas .
Detta är särskilt viktigt för att höja effektiviteten av de beviljade anslagen .
Problem uppstår dock särskilt i och med att anslagen beviljas årsvis och är knutna till projekt , exempelvis Phare , i jämförelse med den flerårsbasis som gäller för Interreg-anslag och det åtgärdsrelaterade anslagsbeviljandet .
Detta kommer framdeles att medföra praktiska problem , men jag hoppas att det ändå blir möjligt att genomföra Interreg på ett meningsfullt sätt .
Herr talman , mina damer och herrar !
Gemenskapsinitiativet Leader har visat sig vara ett verktyg för att ge impulser till innovativ utveckling och till pilotprojekt i liksom från landsbygdsområdet .
Därför är upprätthållandet av just detta gemenskapsinitiativ och den nya upplagan i Leader + -programmet mycket välkomna .
Det nya Leader + -programmet kan nu tillämpas på hela landsbygdsområdet i Europeiska unionen , vilket leder till bättre möjligheter för de projekt som skall stödjas .
Det är viktigt att samordna Leader + med övriga stödmöjligheter i Europeiska unionen , men precis lika viktigt är det att samordna det med de andra nationella stöden .
Det måste undvikas att stöden överlappar varandra , och samtidigt måste synergieffekter kunna utnyttjas .
I enlighet med detta måste målet att stärka integreringen av de olika Leader-stödområdena verkligen välkomnas .
Jordbruket är en av de bärande pelarna på landsbygdsområdet och måste kunna få del i Leader-initiativet , eller också kan den strukturella förändringen i jordbruket få sällskap av Leader-initiativet genom att nya arbetstillfällen skapas på landsbygden .
Alla ekonomiska sammanhang som rör landsbruket måste uppmärksammas i Leader + -programmet , och endast genom gemensamma ansträngningar kan man då nå det optimala .
Leader måste nu förverkligas .
De operativa programmen måste beviljas av kommissionen så snart som möjligt , dvs. en praktiskt genomförd och effektiv hantering av förslagsställandet samt snabbast möjliga godkännande av förslaget .
Fem månader har man räknat med .
Det tycker jag är litet för lång tid .
Man bör i detta fall försöka klara sig med kortare tidsfrister .
För den som har utvecklat ett projekt och fått det färdigt vill också sätta igång med genomförandet så snart det bara går .
Trots all glädje över den nya utformningen av gemenskapsinitiativet Leader + är det dock en sak som ligger mig varmt om hjärtat : Europeiska kommissionen har i sitt förslag krävt ett övervakningscentrum för Leader + -programmet utan att närmare gå in på hur förslaget skall genomföras .
Detta innebär följande frågor för mig : Vem skall arbeta där ?
Hur väljs dessa personer ut ?
Framför allt , varifrån kommer det kapital som behövs , och var skall detta övervakningscentrum vara beläget ?
Jag menar nu att Leader + -programmet inte behöver ett öre till ytterligare förvaltningsuppdrag , vilka det av naturliga skäl i alla fall skulle åligga kommissionen att utföra .
Dessutom visar erfarenheten från andra områden där övervakningscentrer har inrättats att dessa förutom ett tvivelaktig skapande av nya arbetsplatser inte gör någon större nytta .
Jag uppmanar därför kommissionen att själva och direkt sköta sina kontrolluppdrag samt att arbeta för en god utveckling av Leader + -programmen .
Dit hör ju också utvärderingen och offentliggörandet , vilket hittills ju också har varit fallet .
Herr talman !
Den största delen av de gränser som under sekler delat Europa är tillskapade på ett konstlat sätt .
De separerade unika geografiska områden och skapade starka skillnader i form av balanserad utveckling och sammanhållning .
Våra inre gränser , eller det som är kvar av dem , ger inte längre upphov till krig , men de fortsätter att ge upphov till ekonomiska skillnader , sociala gränser och kulturell avskärmning mellan Europas folk .
Från gemenskapens institutioner måste vi arbeta för att komma över denna ärrbildning i gränsområdena , som är en motsättning till andan av europeisk enhet .
Den ekonomiska och sociala sammanhållning som vi kämpar för konkretiseras genom Interreg-initiativet , i den territoriella sammanhållningen och i integrationen av gränsområden och vår kontinents randområden .
Interreg är sedan sin tillblivelse fröet till en verklig gemenskapspolitik för den fysiska planeringen av territoriet och en verklig polycentrisk uppfattning om det europeiska territoriet .
Europaparlamentet beklagar bara att vi måste anta en resolution om detta initiativ , som vi håller med om , när vi ännu inte känner till utvärderingen av Interreg II .
Men vi är medvetna om att det inte är lämpligt att dröja längre med tillämpningen av denna tredje utgåva , eftersom vi då skulle kunna riskera flera projekts framgång och en kontinuitet i de projekt som redan är igång .
Interregs framgångar är uppenbara och det uttrycker de lokala , regionala och nationella myndigheter som deltagit i medfinansierade projekt .
Att lära tillsammans , förnya , dela projekt och goda erfarenheter , förstå och tolerera varandra är några av de lektioner som deltagarna i detta initiativ kan lära av detsamma .
Det finns en hel del intressanta frågor kring detta , observation , koncentrationsprincipen ...
Jag skulle vilja uppehålla mig kring de förvaltande organen .
Det är nödvändigt att söka gemensamma , interregionala och transnationella förvaltningsorgan i vilka alla lokala och regionala myndigheter deltar aktivt , samt de ekonomiska och sociala parterna .
Parallella projekt på ena och andra sidan gränsen bör inte upprepas .
Vi måste skapa en gränsöverskridande kultur och för detta ändamål är det nödvändigt att finna nya vägar när det gäller administrativt samarbete och med fantasi övervinna existerande hinder , samt övervinna de svårigheter de olika graderna av kompetens i varje medlemsstat , i varje region och i varje kommun innebär .
Det får inte vara så att ett projekt inte kan genomföras på grund av samtalssvårigheter .
Under diskussionerna i utskottet har vi också konstaterat svårigheten att samordna Interreg med andra finansiella instrument av årlig eller tvåårig karaktär , som Meda , Tacis eller Phare .
Genom förslaget till resolution i parlamentet har man verkligen försökt uppmärksamma dessa svårigheter genom att formulera förslag till kommissionen som gör det möjligt att lösa dem och genom att uppställa rimliga tidsfrister för att genomföra nödvändiga ändringar .
Herr talman !
Mitt skäl till att bidra till denna debatt har att göra med att Urban-initiativet - särskilt i Irland - har varit mycket framgångsrikt och jag vill verkligen att Europeiska unionen ger ytterligare bidrag på detta område .
Det är ett tråkigt faktum att det finns flera hundra , om inte tusentals , samhällen i Europeiska unionen som lider av en mycket allvarlig fattigdom och eftersatthet .
T.o.m. i medlemsstater och städer som är oerhört välmående finns det många som bor i getton , under levnadsbetingelser där det inte finns tillräckligt med moderna bekvämligheter , där utbildningen är bristfällig , där den fysiska infrastrukturen är underutvecklad och där narkotika och andra fenomen är mycket vanliga .
Det verkar som om Europeiska unionen , för att visa att den har en roll när det gäller att hjälpa Europeiska unionens medborgare , måste hjälpa medlemsstaterna för att visa att unionen fungerar för dessa medborgare och deras familjer .
Programmet har varit oerhört framgångsrikt i Irland , på samma sätt som jag naturligtvis känner till att det varit framgångsrikt i andra länder .
Det var litet långsamt under inledningsfasen här , men detta berodde på att det var nödvändigt att lokalbefolkningen själv utvecklade dessa program .
Det är viktigt att de använder sin initiativkraft och sin egen kännedom om lokala förhållanden vid utvecklingen av detta initiativ .
Det skulle vara mycket lätt att se till att få dessa program snabbt utvecklade och i rätt tid om man tog hjälp av externa sakkunniga , men detta skulle undergräva hela syftet med Urban-programmet .
Jag vill ta upp ytterligare en sak innan jag slutar : vi bör ställa krav på det sätt på vilket dessa medel tilldelas och den plats detta program utvecklas , i det avseendet att det sker i samband med en seriös Urban-utvecklingspolitik .
Detta är tyvärr inte fallet i Irland .
Jag applåderar det innovativa förhållningssättet inom Equal-programmet och målet att få ut diskriminerade grupper på arbetsmarknaden .
Utvecklingspartnerskapen är en mycket klok idé , trots att de befinner sig på experimentstadiet .
Det finns emellertid framför allt två skäl till varför jag har betänkligheter rörande utvecklingspartnerskapen .
De borde vara tillgängliga för mindre grupper , tillgängliga i det avseendet att de skall kunna planera , genomföra och övervaka programmen .
Vi måste ha ett stort mått av flexibilitet inom programmet .
Jag har också innan uttryckt oro rörande användningen av jargong i stället för ett enkelt och tydligt språk , så att det blir tillgängligt för alla .
Jag är glad att denna tanke godtogs i betänkandet , men jag kan inte stödja ändringsförslag 9 , eftersom detta ändringsförslag faktiskt inte alls skrivits på ett enkelt språk .
För det andra oroar det mig att vissa diskriminerade grupper har särskilda problem - t.ex. de handikappades situation i fråga om tillträde till sina arbetsplatser .
Genom projekten bör man också särskilt ta itu med detta problem .
Man bör titta på dessa frågor samtidigt som man fastställer programmen .
Jag har sannerligen för avsikt att göra detta tillsammans med organisationer och grupper i min valkrets i West Midlands .
Låt mig nu ta upp den kontroversiella frågan om asylsökande och flyktingar .
Även om jag inte stöder att de flyktingar som förvägrats flyktingstatus och hotats med avvisning skall få tillgång till Equal-initiativet , stöder jag möjligheten till tillgång för alla övriga asylsökande och flyktingar .
Det är bara rätt och riktigt att de skall kunna få tillgång till Equal-initiativet på samma sätt som alla andra .
Herr talman , kära kolleger !
I betänkandet om Leader är det landsbygdens utveckling som står i centrum .
Det är inte så vanligt och det är därför glädjande , särskilt som Leader-programmen varit huvudbeståndsdelar i unionens politik för landsbygdsutveckling .
Det bör erinras om att dessa program inte bara varit strukturerande beståndsdelar för en politik för fysisk planering utan också grundläggande instrument för ekonomisk och social sammanhållning i områden som ofta är ömtåliga , exempelvis områden med utbredning av ödemark .
Det är viktigt att betona att för att kunna komma i fråga för stöd enligt Leader-programmet har de lokala aktörerna samarbetat , diskuterat och utarbetat projekt .
Därför har dessa program varit viktiga för en demokrati där människor är delaktiga och för medborgartanken i Europa .
Konceptet Leader + skall också innehålla alla positiva aspekter av tidigare program .
En viktig fråga uppstår alltså : varför skall vi efter att i tio år framgångsrikt ha bedrivit dessa program förpassa Leader + till en experimentroll ?
Finns det så många andra europeiska åtgärder som gör att man kan stoltsera med 800 originella specifika erfarenheter som varit ovanligt lyckade ?
Hur länge tänker kommissionen fortsätta att behålla Leader på experimentstadiet innan programmet tillåts ingå i det allmänna konceptet för landsbygdsutvecklingens mainstreaming ?
Jag ställer mig också frågande till de minskade riktlinjer dit kommissionen vill förpassa Leader + .
Herr kommissionär !
När vi européer , efter Seattle , kämpar för de många funktionerna i projekten för landsbygdsutveckling , varför då begränsas av kriterier med mycket otillräckliga medel ?
Det är en miljöpartist som talar till er : försiktighetsprincipen och en hållbar utveckling kräver ett mycket mer varierat synsätt under många fler former .
I det sammanhanget föreslår kommissionen att vi ytterligare skall begränsa åtgärderna för samarbete med lokala aktionsgrupper till enbart kandidatländerna .
Det skulle vara bättre , vilket också utskottet för regionalpolitik föreslår , att ha en förstärkt samordning mellan Leader + och gemenskapens program för samarbete och partnerskap , såsom Interreg , Phare , Sapard eller Meda .
Att vara solidarisk med Östeuropa är nog bra , men det räcker inte .
Traditionen från de tidigare programmen , med länderna i söder , särskilt kring Medelhavet , får inte överges .
Därför kan vi ännu en gång betona att det som saknas på jordbruksområdet och inom landsbygdsutvecklingen är medbeslutande , som skulle göra det möjligt för oss att verkligen få medel för att program som kräver samarbete och tvärgående åtgärder skulle kunna innebära framsteg .
Herr talman !
Jag har några mycket korta kommentarer .
Vi diskuterar den nya programplaneringsperioden och de nya riktlinjerna för de fyra gemenskapsinitiativen , utan att ha tillgång till en egentlig och fullständig utvärdering av den föregående perioden .
Det är mycket negativt .
Programmen och målen är vanligtvis väldigt optimistiska , resultaten är emellertid inte alltid tillfredsställande , och ofta lämnar bristen på öppenhet i förening med projektens komplexitet stort utrymme för misshushållning och till och med bedrägerier .
De gemenskapsinitiativ som vi diskuterar kan under vissa omständigheter spela en positiv roll .
Det är dock nödvändigt att de inte underställs mål och strävanden inom ramen för en mer allmänt negativ ekonomisk och social politik , utan att de utvecklar en egen , självständig roll .
Till exempel innebär Equal-initiativets anpassning till målen om anställbarhet och ökad elasticitet i förhållandet mellan arbetsmarknadens parter att det förvandlas till en ny version av de lokala sysselsättningspakterna .
Utvidgningen av Leader-initiativet till alla unionens områden innebär en risk för en ytterligare marginalisering av de mindre gynnade regionerna , till fördel för de mer utvecklade regionerna .
Interreg-initiativet skall omfatta utvalda regioner , med särskilt betoning på randregioner , öregioner , bergs- och icke-bergsregioner , som till exempel Artas län i Grekland , som helt felaktigt har utelämnas i bilaga I till kommissionens meddelande .
Herr talman !
Detta parlament och kommissionen har bestämt att landsbygdsutveckling skall betraktas som ett prioriterat politikområde , och jag vill här i dag välkomna den ansvarige kommissionären , kommissionär Fischler .
Vår reaktion i samband med de stödbehov som finns på landsbygden har varit långsam , men jag antar att det är bättre sent än aldrig .
Familjejordbruket har nu erkänts som ett viktigt inslag i den europeiska jordbruksmodellen och är ett mål som skall diskuteras inom ramen för Agenda 2000 .
Jag anser att det inom de kommande fem åren kommer att fattas beslut som bestämmer framtiden för tusentals familjejordbruk som befinner sig på marginalen .
Det anstår oss alla att göra allt som står i vår makt för att säkerställa deras fortlevnad .
Som kommissionären känner till kommer inte bara jordbruksnäringen att vara tillräcklig för att säkerställa en hållbar utveckling på landsbygden .
Av detta skäl behöver vi en samordning av alla politikområden som kan spela en positiv roll för landsbygdens utveckling .
I detta avseende har Leader etablerats som ett effektivt utvecklingsinitiativ .
Det ger möjligheter för lokala samhällen att fastställa sin utvecklingspotential och att aktivt delta i en diskussion av dessa problem .
Det frivilliga deltagandet i utvecklingsprogram är inte alltid något som uppskattas fullt ut .
Genom Leader kan det emellertid inte råda några tvivel rörande effektiviteten i detta sammanhang som en integrerad del av en bredare EU- och nationell politik .
Samtidigt som jag sammanfattningsvis välkomnar godkännandet av Leader + , oroas jag av tidsglappet mellan avslutandet av Leader II och inledningen av det nya programmet .
Jag uppmanar er att ta allvarligt på detta problem .
Ett avbrott i verksamheten kommer att få allvarliga konsekvenser för programmet och en störande effekt på de frivilliga och yrkesmässiga arbetsinsatserna .
Herr talman , herr kommissionär , mina damer och herrar !
Efter att ha fått kännedom om meddelandet från kommissionen om initiativet Interreg III , och med tanke på att jag inom ramen för utskottet för regionalpolitik , transport och turism deltagit i omröstningen om Decourrières betänkande , vill jag inte bara uttryckligen säga att vi principiellt är överens dels om initiativet , såsom det föreligger , och särskilt inom ramen för Interreg III B , och dels om att kommissionen skall godkänna den verksamhet som bidrar till att återupprätta landskap som lidit skada på grund av jordbrukspriserna , en sektor där ett stort antal föreningar , särskilt på jaktområdet , redan gör enorma satsningar i mitt land .
Jag vill också ge mitt uttryckliga stöd till kommentarerna från utskottet för regionalpolitik , transport och turism , framför allt när det gäller att beklaga bristen på integration av de yttersta randområdena inom område A i programmet , eller påpeka bristen på precision när det gäller urvalskriterierna för villkoren för genomförande av område III C , och slutligen när det gäller att kräva att parlamentsledamöterna skall vara delaktiga i ett europeiskt övervakningscentrum för gränsöverskridande , transnationellt och interregionalt samarbete .
Jag vill också uttrycka ett verkligt förbehåll mot tendensen i kommissionens meddelande att , enligt Interreg III och III B , knyta miljöskyddet enbart till utvecklingen av Natura 2000 , som förefaller mig ofta vara ett alltför abstrakt medel för att försvara de ekologiska system , vars användare riskerar att uteslutas eller starkt begränsas .
Jag skulle avslutningsvis vilja betona , genom att i förväg be om förståelse från kommissionen och berörda ministerråd , att det skulle vara lämpligt att ytterligare informera de europeiska folkvalda om de förfaranden som är knutna till inrättandet av Interreg-ärendena och liknande initiativ .
Och vi måste dessutom ytterligare införliva dem i processen med att utarbeta och genomföra berörda program , annars blir det svårt att förstå och försvara deras roll mot lokala och nationella myndigheter och till och med mot medborgarna .
Herr talman !
Först och främst skulle jag vilja framföra ett hjärtligt tack till föredraganden för Equal-betänkandet , Stenzel , för allt som hon har gjort för att för att vi allesammans skall få insikt i detta svåra ärende .
Equal är ett mycket svårt program eftersom man där försöker att sammanföra så många gamla program och ändå vill se över dem på ett nytt sätt , och detta med mindre pengar än vad som stod till förfogande i de tidigare fonderna .
Det är en svår uppgift .
Det är bara antalet personer som berörs av dessa program som egentligen inte har minskat .
Därför är det mycket svårt att få en balans till stånd , inte bara mellan de olika länderna , inte bara mellan de olika delarna , utan i synnerhet även mellan de olika grupper som nämns i programmet , och det är egentligen det som har sysselsatt oss fram till i dag .
Här och där fälls kommentarer om att den ena gruppen måste få mer än den andra .
Själv har jag särskilt ägnat mig åt de handikappades och de äldres ställning inom ramen för programmet , och jag måste säga att de handikappade och de äldre hade kunnat bli helt bortglömda om inte Europaparlamentet hade ägnat sig åt den frågan så intensivt .
En del andra grupper har nämnts , men det är framför allt medlemsstaterna som ligger på lur .
Jag känner till exempel till en medlemsstat som vill använda en stor del av hela programmet till en enda del , nämligen flyktingarna .
Jag skulle därför vilja be kommissionären att ordentligt se till att det upprättas en balans mellan de olika grupperna .
Det får inte vara så att en medlemsstat , genom att åberopa subsidiaritetsprincipen som förevändning , kan säga att allt skall gå till en enda grupp .
Jag tror att det krävs sträng tillsyn i detta fall , för annars får man just det som Meijer varnade så starkt för , nämligen att det kommer att uppstå etablerade intressen och att människor tänker att pengarna är deras .
Det är inte på det sättet !
De måste varje gång fördelas på nytt .
Det skall handla om innovativa projekt , och det får inte vara så att de helt och hållet försvinner in i finansministerns kassa .
Det är inte syftet , och det är en viktig punkt som vi måste beakta här .
Jag tror att de kvarvarande problem som vi har haft inom parlamentet , som till en stor del härstammar från det faktum att det är så svårt att göra denna avvägning , kan lösas .
Vad kommissionen beträffar hoppas jag att den kommer att kunna ansluta sig till den kompromiss som kommer att nås här i parlamentet och som framför allt är inriktad på balans .
För att ytterligare understryka detta - situationen är naturligtvis aningen svår - har parlamentet för enkelhetens skull och för säkerhets skull tills vidare placerat Equal-programmet i reserven , så att parlamentet så småningom skall bli övertygat om på vilket sätt genomförandet kan komma till stånd .
Jag tror att det också är positivt .
Parlamentets ställning i hela denna procedur är litet otydlig .
Även i arbetsordningen är denna ställning otydlig , och just därför är det mycket bra med denna reserv .
Herr talman !
Värderade kolleger !
Det är ett oemotsägligt faktum att Interreg-initiativet stöder ansträngningarna att nå ekonomisk och social sammanhållning i Europeiska unionen .
Jag vill dock betona den särskilda betydelse som Interreg har för Balkanregionen , där de senaste årens politiska utveckling och krigshandlingar har fått stora ekonomiska konsekvenser för grannländerna , särskilt för mitt land , Grekland , som är det enda medlemslandet som är beläget på den hårt drabbade halvön .
För Grekland , grannländerna Italien och Österrike , men även för hela Europa , är Balkans sociala och ekonomiska återuppbyggnad , som skall leda till politisk stabilitet , en fråga av största betydelse .
Fram till i dag har vissa av länderna på Balkan fått stöd genom Phare- och Obnova-programmen , andra inte .
Under den nya programplaneringsperioden , inför utvidgningen och med hänsyn tagen till att stöd genom nya stödinstrument och förordningar , som till exempel Ispa och Sapard har planerats , är det absolut nödvändigt att samordna stödet på Interregs tre insatsområden med det övriga stödet till tredje land .
Vi välkomnar följaktligen formuleringarna om detta i kapitel 7 i Europeiska unionens text om fastställande av Interreg-riktlinjer .
Ansträngningarna för att samordna och följaktligen effektivisera planeringen måste fördelas lika på alla program , och jag säger detta eftersom det i Meda-programmet , under den föregående perioden , fanns vissa problem som bör lösas , så att vi behandlar alla de tredje länder som deltar i programmet lika .
Jag skulle vilja avsluta , herr talman , med att konstatera att man i den nya planeringen av områdena för mellanstatligt samarbete inte har tagit hänsyn till Medelhavsområdets geografiska egenhet , som borde rättfärdiga skapandet av ett särskilt område för kust- och öregioner .
Vi begär alltså av kommissionen att den särskilt skall beakta frågan om samarbete i havsnära regioner och i öregioner vid kommande revideringar av områdesplaneringen .
Avslutningsvis , herr talman , betonar jag nödvändigheten av att Europeiska unionen insisterar på denna slags initiativ , som avser att utplåna orättvisor mellan våra regioner och att få till stånd en harmonisk utveckling för dem .
Och eftersom det i dag är Alla hjärtans dag , föreslår jag , som gammal borgmästare i en regional stad , att vi alla förklarar vår kärlek till de europeiska regionerna , de som behöver den kärleken .
Herr talman , bäste kommissionär Fischler !
Vid utvecklingen av landsbygden kan och måste man ta hänsyn till tre problemställningar , nämligen bibehållandet av sysselsättningstillfällen , landskapsvården och inte minst den lokala kulturen , för den är viktig !
Endast om befolkningen kan stanna kvar på landet kan livskvalitén på landet förbli garanterad på sikt .
Vad flykten från landsbygden innebär kan vi iaktta i vissa områden i Alperna , och följderna är katastrofala !
Men jag vill varna för att med detta program överföra stadskulturen till landsbygden .
Och vi skall heller inte skapa bidragsberoende strukturer som för all framtid blir hänvisade till stöd .
För att trygga en hållbar utveckling - ett slagord som med tiden blivit ganska tomt , men vi alla förstår vad vi menar med det - krävs det bland annat att turism och jordbruk integreras på landet .
Investeringarna måste gå i en visionär riktning .
Unga kreativa individer måste kunna hållas kvar på landsbygden .
Om de allihop flyttar händer det inte så mycket mer där .
Ingen av oss är särskilt förtjust i principen om att alla ges lika mycket oavsett behov , och projekten av pilotkaraktär måste så att säga dra med sig andra liknande projekt som en lavin .
Jag pläderar för att slutna kretslopp skall stödjas , och även om Leader II och Leader II här och där har haft sina brister så var resultatet säkerligen positivt ändå .
Jag vill be alla fundera över att inte bara bevilja undantag i nordliga länder , utan även för bergsområdena , Alperna , Pyrenéerna , Sierra Nevada som jag just kommer ifrån , nämligen i fråga om invånarantal och befolkningstäthet .
( Applåder ) Herr talman !
Jag vill tala om Equal-betänkandet , särskilt frågan om flyktingpolitik .
I förra veckan diskuterade vi den österrikiska regeringsbildningen med stort engagemang .
I dag diskuterar vi redan den österrikiska regeringskoalitionens flyktingpolitik , eftersom Stenzel som har författat Equal-betänkandet ju representerar det österrikiska konservativa regeringspartiet och dess politik .
Det mest uppseendeväckande i hennes ursprungliga betänkande var att hon ville begränsa flyktingstödet till den lilla grupp flyktingar som omfattas av Genèvekonventionen , dvs. så kallade kvotflyktingar eller FN-flyktingar .
I själva verket är det de andra flyktingarna , nämligen de som står utanför kvoten och FN-stöd , som har det största behovet av stöd .
Utskottet förkastade detta diskrimineringsförslag och beslutade att alla flyktingar skall få plats i Equal-programmet på lika villkor .
En del av utskottet solidariserade sig emellertid med Stenzels förslag och formuleringar .
Det betyder enligt mitt sätt att se att Haiderpolitiken redan kastar sin skugga över detta parlament .
Därför är det av avgörande betydelse att kammaren med största möjliga eftertryck slår fast att alla flyktingar skall ha plats i Equal-programmet .
Jag vill till sist säga att jag hade vissa betänkligheter i förra veckan när vi diskuterade regeringsbildningen , men när det gäller att diskutera och kritisera den österrikiska flyktingpolitiken , då har jag inga betänkligheter .
Jag hoppas att engagemanget i kammaren blir lika stort denna gång .
Herr talman !
Under EU : s senaste budgetplan från 1994 till 1999 , när det fanns 13 olika initiativ i kraft , var det gränsöverskridande Interreg II-programmet ett viktigt initiativ .
Det faktum att nästa strukturfondsrunda mellan 2000 och 2006 omfattar Interreg-initiativet anser jag vara en mycket tydlig fingervisning om den betydelse som tillmäts detta av EU : s medlemsstater .
Interreg I-programmet mellan 1989 och 1993 och Interreg II-programmet mellan 1994 och 1999 har visat sig vara en fullständig framgång när det gällt att skapa ett närmare samarbete mellan angränsande medlemsstater i frågor som rör social och ekonomisk utveckling .
Eftersom jag själv kommer från gränstrakterna i nordvästra Irland har jag sett den viktiga roll som Interreg I och II har spelat under årens lopp , och jag är glad att kunna välkomna Interreg III .
Kommissionen kommer att tilldela 67 miljoner pund till Interreg III-programmet , som kommer att användas till en fortsatt utveckling av gränsöverskridande ekonomiska projekt mellan Irland och Nordirland .
Europeiska unionen har spelat en viktig roll vid utvecklandet av gränsregionerna i Irland under årens lopp .
Europeiska unionen är den enskilt största bidragsgivaren med 80 miljoner pund till Internationella fonden för Irland .
Europeiska unionen bidrar med 75 procent av det totala Freds- och försoningsprogrammet .
Sammanfattningsvis har Interreg , Internationella fonden för Irland och Freds- och försoningsprogrammet spelat en viktig roll för den löpande fredsprocessen .
Herr talman !
Jag skall tala om Interreg och bland annat för att respektera tidsbegränsningen hålla mig till några få kritiska punkter .
Vi har alla gett uttryck för en positiv syn på att detta program förlängs och på utvidgningen av insatsområdena till att förutom samarbete över gränserna även omfatta samarbete mellan nationer och regioner .
Detta hindrar dock inte att vi är medvetna om det faktum att större delen av resurserna - mellan 50 och 80 procent - kommer att reserveras för samarbetet över gränserna , för volet A i Interreg III-programmet .
Det val man sedan har gjort , att för detta volet befästa de nuvarande samarbetsområdena , vad gäller vilka regioner som äger tillträde , anser vi fortfarande är både felaktigt och motsägelsefullt .
Vi hoppas verkligen att kommissionen kommer att se över detta och vidgå parlamentets ståndpunkt i sak , och inte som en formell aktningsbetygelse .
Samarbetet över gränserna sker fortfarande nästan uteslutande över landgränserna och på de ställen man har gjort undantag för vattengränser saknas insyn i besluten och de bär ofta spår av kompensation för andra delar av gemenskapspolitiken .
Diskrimineringen framstår som enormt mycket allvarligare för öarna , vilkas regionala förhållanden inte kan annat än präglas av att de uteslutande har havsgränser .
Detta är i linje med en diskriminering som man fortsätter att tillämpa utan att ta hänsyn till artikel 158 i fördraget , som gäller öregionerna i sammanhållningspolitiken .
Det är ännu mer allvarligt att detta sker utan hänsyn till den nya väg vi har slagit in på i och med utvidgningen till regioner som Malta .
Härav de förslag vi har lagt att utvidga de regioner som kan komma i fråga åtminstone till Siciliens Nuts III-gränser gentemot Malta och för alla de adriatiska regionerna gentemot Balkan .
Herr talman , herr kommissionär , kära kolleger !
Jag skulle vilja uttrycka min tacksamhet över att kunna konstatera att de yttersta randområdena , däribland de franska utomeuropeiska departementen , varit föremål för ett visst intresse inom ramen för initiativet Interreg III , vilket öppnar nya perspektiv för att de skall kunna samarbeta med länderna inom sitt geografiska område , även om man kunde ha hoppats på något bättre , bl a när det gäller tillgång till de olika områdena .
Under lång tid har våra regioner haft blicken fästad på sin europeiska huvudstad , sannolikt en kvarleva från kolonialtiden , och struntat i och till och med föraktat sina närmaste grannar .
Detta hör i dag absolut till det förgångna .
Våra regioner har blivit medvetna om att de tillhör en miljö som de är knutna till , inte bara geografiskt utan också genom sin kultur och sitt folks historia , vilket ger upphov till en stark strävan efter en djupare förankring i denna miljö .
Men denna insikt handlar inte bara om identitet .
Den är också beroende av en rättvis uppskattning av våra tillgångar .
La Réunion befinner sig exempelvis mitt i axeln för utbyte mellan länderna i södra Afrika och de i Sydostasien .
Ön kan inte stå vid sidan om de regionala grupperingar som verkar i området , eftersom den då riskerar att gå miste om en historisk möjlighet , och detsamma gäller våra regioner i Västindien .
Avslutningsvis är vi övertygade om att våra ungdomar kan skönja en utväg ur den dramatiska arbetslösheten som gör dem förtvivlade , om vi till intilliggande länder kan exportera den know-how som förvärvas tack vare strukturfondernas åtgärder .
Utnyttjandet av Interregs anslag kan göra våra regioner till verkliga brohuvuden för Europeiska unionen inom deras geografiska områden , och på så sätt ge dem en världsomspännande dimension .
Jag räknar med kommissionen och särskilt med er , herr kommissionär , för att ge dem medel till effektiva åtgärder .
Herr talman , kommissionärer !
Jag välkomnar varmt möjligheterna till ett ökat europeiskt samarbete i samband med Interreg , men jag oroar mig för att förslaget ger färre möjligheter för havsområdena än för andra områden i detta avseende .
Jag förstår kommissionens egen oro över att geografiskt avstånd kan inverka menligt på ett effektivt samarbete .
Det finns i vilket fall många havsområden som redan upprättat kontakter .
Olika lokala myndigheter i Nordsjöområdet är ett bra exempel på detta .
Interreg skulle mycket väl kunna förstärka detta samarbete .
Som ett resultat av detta vill jag se att det görs vissa mindre ändringar av riktlinjerna för att skapa litet mer flexibilitet och för att anpassa de sätt på vilka havsområdenas intressen kan hamna mellan område A och område B. Dessa anpassningar omfattar ett förtydligande av möjligheterna för samarbete mellan havsområden och tillåtande av en bredare utveckling av praktiska och genomförbara projekt , i synnerhet de som har en infrastrukturell karaktär .
Sådana åtgärder kommer att likställa havs- och öområden med andra områden i EU .
Jag hoppas att de blir antagna .
Herr talman !
Vår grupp välkomnar den övergripande kraften hos Equal-initiativet genom att , om du är en brittisk muslim som har någon form av fysiskt handikapp inte längre behöver välja mellan vilken diskrimineringskategori man tillhör som målgrupp : Man kan använda sin sakkunskap och erfarenhet för att lösa problem , i stället för att betraktas som själva problemet .
Det finns mycket sakkunskap inom de relevanta organisationerna som är värd att dela med sig av .
Vi välkomnar också erkännandet av behovet av utvärdering och spridning av bästa metoder för åtstramning av den gränsöverskridande nivån .
Vi är därför bekymrade över , som andra har nämnt , antalet ändringsförslag som försöker att ytterligare marginalisera en del av de i samhället som redan tillhör de mest marginaliserade , genom att förespråka en mycket snäv definition av " flykting " .
Min grupp kommer inte att stödja dessa ändringsförslag .
Vi är också bekymrade över det antal ändringsförslag som innebär att man genom att försöka införa en större flexibilitet , kanske löper en risk att skapa förvirring när det gäller var ansvaret för Equal-initiativets verksamhet ligger .
Herr talman !
Det gläder mig att se att Urban-initiativet ges en mer helhetlig inriktning och att man med initiativet försöker lösa sammanhängande problem .
Det finns dock , herr talman , en risk med denna utspridning : att våra försök att uppfylla många mål leder till en övergripande ineffektivitet .
Varje enskilt fall av tillbakagång i ett stadsområde är naturligtvis speciellt .
Det finns emellertid en resultant , en hård kärna , som består i att arbetslösheten ökar , att de offentliga tjänsterna försvinner eller skärs ned samt att små och medelstora företag , affärer och andra inrättningar försvinner .
Jag skulle önska att man med Urban-initiativet först och främst riktade in sig på att försöka finna svar på dessa orsaker till tillbakagång i städerna .
Och då är det naturligtvis nödvändigt att nå samförstånd och att samordna den centrala politiken med utvecklingspolitiken , så att även denna ges en ny inriktning och samverkar med målen i de Urban-initiativ som genomförs i våra länder , i stället för att helt enkelt lägga fram de där programmen som ett alibi för frånvaron av en sådan politik .
Herr talman , herr kommissionär , kära kolleger !
Jag begränsar mitt inlägg till Francis Decourrières betänkande .
Programmet för gemenskapsinitiativet Interreg är ett extremt viktigt verktyg när det gäller europeisk utveckling och fysisk planering , särskilt om vi effektivt skall beakta förhållandet mellan Europeiska unionens centrum och dess randområden .
Interreg skall därför vara ett instrument som främjar unionens territoriella sammanhållning , om vi vill undvika ett europeiskt territorium uppdelat i två eller tre hastigheter .
Det förefaller mig självklart att de regionala och lokala myndigheterna , de organisationer som företräder dem , Regionkommittén och självfallet Europaparlamentet , tydligare och så snart som möjligt skulle ha kopplats in när det gäller att utarbeta programmet .
Men man måste konstatera att så inte var fallet när kommissionen förberedde sitt meddelande , som offentliggjordes den 13 oktober förra året .
Även om jag godkänner de allmänna riktlinjerna för Interreg III , förefaller det mig ytterligt viktigt att se till att det finns en bättre förbindelse mellan detta program - som finansieras av Europeiska regionala utvecklingsfonden ( ERUF ) - och övriga fonder för yttre samarbete , däribland bl.a.
Europeiska utvecklingsfonden avsedd för AVS-länderna .
I det hänseendet skulle jag vilja tacka utskottet för regionalpolitik , transport och turism för att ha antagit ett av mina ändringsförslag som lägger till Europeiska utvecklingsfonden ( EUF ) i förteckningen över dessa fonder .
De yttersta randområdena , bl a de fyra franska utomeuropeiska departementen , måste kunna samordna Interreg III och EUF för att också de skall kunna finansiera samarbetsprojekt med sina AVS-grannar inom respektive geografiska område .
Jag ber också kommissionen att vänligen på nytt överväga de dåliga möjligheter som erbjudits de yttersta randområdena och öregionerna enligt riktlinjerna i meddelandet .
Dessa regioner skall , liksom samtliga övriga regioner i unionen , kunna utnyttja Interreg III fullt ut , särskilt som programmet Regis , som var avsett för dem , nu avskaffats .
Avslutningsvis vill jag beklaga de låga ekonomiska bidrag som avsatts för område C , avsett för samarbete mellan regioner , och vars betydelse inom gemenskapen ändå inte kan förnekas .
Herr talman !
Min utgångspunkt är Equal-betänkandet och jämställdhet mellan män och kvinnor , även om jag måste erkänna att det emellanåt är tröttsamt att tala om denna fråga som har fått upprepandets natur , i varje fall när man är i min ålder .
Men det är tyvärr nödvändigt att återigen påpeka att vi inte uppnått jämställdhet .
Men kanske kan ett genombrott här leda fram till ändringar på andra områden .
För mig betyder nämligen inte jämställdhet att båda parter i ett äktenskap arbetar hela tiden och lämnar barnen till en dagmamma , dvs. en invandrare , som inte har fått en chans att få ett annat jobb .
Om det skall vara så har vi inte kommit någonvart sedan solkungarnas tid .
Nej , jämställdhet innebär att vi alla deltar i både arbetslivet och familjelivet .
Utvecklingen går tyvärr inte i den riktningen , tvärtom .
Jag tycker därför att punkt 7 innehåller något mycket viktigt .
Här står nämligen : " Equal kommer att användas som försökslaboratorium för utveckling och förmedling av nya metoder för genomförande av sysselsättningspolitik " .
Man får hoppas att det lyckas .
Herr talman !
I samband med arbetsordningen vill jag bara säga att om jag inte är här när kommissionen svarar - inte därför att jag ställt några särskilda frågor , men jag hoppas dock att kommissionen har gjort efterforskningar - beror detta på att det samtidigt med denna debatt pågår ett sammanträde i utskottet för kvinnors rättigheter och jämställdhetsfrågor om kvinnor i beslutsprocessen .
Herr talman , mina damer och herrar !
De som ägnar sig åt landsbygdsområdet vet att Leader-programmet , såväl Leader I som Leader II - och jag hoppas även Leader + - hör till berättelserna om de framgångar som Europeiska unionen har lanserat .
Framgångarna kom sig även av att Leader-programmens grundkoncept framkallade en mycket stor aktivitet hos den berörda befolkningen .
Det gläder mig att grundsatsen för Leader + har stannat vid detta grundkoncept .
Det finns dock ett problem som vi måste ta itu med gemensamt .
Eftersom Leader är något som kan liknas vid en verkstad med ett bottom-up-koncept , är det enormt många idéer som under årens lopp har mognat genom Leader I och II , idéer som så småningom förstås inte är så helt nya och framgångsrika längre .
Och på grund av framgångarna leder grundsatsen naturligtvis till att de en vacker dag faller bort ur Leader .
Därför måste vi se till att det som har visat sig vara framstående i de bra Leader-projekten inte plötsligt avbryts , utan de idéer som har visat sig vara goda någon gång måste föras över till de normala programmen som en fast , positiv komponent i stödet till landsbygdsområdet .
Det är ju också grundidén .
Att genom nya idéer i Leader prova något , tillsammans med de inblandade på plats , med de kommunala sammanslutningarna på plats , med många oberoende organisationer , med kyrkorna , tillsammans med alla som har hjälpt till att verkligen få igång nya idéer på landsbygden .
Här måste vi se till att de positiva saker som verkligen sticker ut på något sätt blir en fast beståndsdel i ett förnuftigt arbete inom landsbygdspolitiken .
Nu ber jag kommissionen : Ge akt på att de organisationer och de befolkningsdelar som satsar sin kompetens också verkligen tas emot .
Det får inte vara så att man försöker sig på att mer eller mindre marginalisera den eller den organisationen som bildas just för att bidra med en ny idé och som ännu inte är särskilt känd - och må det så vara på grund av officiell politik på lokal eller regional nivå .
Stanna kvar vid de positiva erfarenheter som Leader hittills har visat .
I början kan det ibland vara litet som att lägga ut rökridåer att säga att det är för idealistiskt uttänkt .
Och sedan under arbetets gång , under genomförandet , framträder det så småningom något som den officiella politiken - även vi på vår nivå - inte alls kunde föreställa sig , att det plötsligt skulle mogna och bli så bra .
Det är detta som har varit charmen med Leader , och det får bara inte gå förlorat !
Herr talman !
Jag välkomnar Equal-initiativet och betänkandet i vilket man betonar behovet av att skilja mellan åtgärder för bekämpning av diskriminering av kvinnor och åtgärder för bekämpning av diskriminering av minoritetsgrupper .
Kvinnor tillhör ingen minoritet och kvinnor drabbas ofta av dubbel diskriminering som medlemmar av minoritetsgrupper , såväl som på grund av sitt kön .
Detta är skälet till varför det behövs särskilda åtgärder för kvinnor , såväl som mainstreaming .
Detta tas upp i betänkandet och man föreslår en integrering av åtgärder för att åstadkomma jämlikhet mellan kvinnor och män i alla arbetsaspekter ; man tar också upp betydelsen av samarbete med de lokala och regionala organ som finns närmast medborgarna , för att se till att alla projektresultat har granskats ur ett jämlikhetsperspektiv .
Deltagandet av frivillig- och gemenskapsgrupper kommer också att bli en viktig del av Equal-initiativet och projekten .
Utvecklingspartnerskapen inom ämnesområdena , vilka anges i ändringsförslag 22 , skulle göra det möjligt även för de mindre organisationerna att spela en roll inom Equal-initiativet .
Min grupp kommer att stödja ändringsförslag 22 .
Herr talman , ledamöter !
Det betänkande kammaren diskuterar i dag är otvivelaktigt mycket viktigt .
Styrkan i gemenskapsinitiativet Interreg för programplaneringsperioden 2000-2006 är , förutom de mål det syftar till , det mervärde det innebär i ljuset av den numera snart förestående utvidgningen av Europeiska unionen till att omfatta nya länder i Östeuropa och Medelhavsområdet .
Det är just inför denna händelse som Europeiska unionen enligt min mening måste ta krafttag för att minska de regionala skillnaderna och sätta stopp för gränsområdenas isolering .
De sistnämnda har faktiskt - det bör man komma ihåg - en viktig roll att spela : rollen som broregioner gentemot de kandidatländer som kommer att bli medlemmar i unionen .
Det är just mot bakgrund av detta som jag har lagt fram några ändringsförslag som jag anser är ytterst viktiga och som utskottet för regionalpolitik , transport och turism har gjort till sina .
Med dessa vill vi utöka de områden som kan komma i fråga för samarbete över gränserna till alla adriatiska regioner liksom de sicilianska provinser som har gräns mot Malta - kandidatland i utvidgningen - vilka i dag oförklarligt nog inte omfattas av avsnitt A i bilaga 1 .
Jag förlitar mig på att kommissionär Barnier och Europeiska kommissionens ordförande tar vederbörlig hänsyn till parlamentets ståndpunkt i frågan , i enlighet med uppförandekoden .
Det är ett grundläggande intresse för hela Europa att främja samarbete med kandidatländerna och ingripa till stöd för gränsregionerna .
Slutligen anser jag att det är önskvärt att man söker förbättra samordningen mellan Interreg-initiativet och de redan befintliga gemenskapsprogrammen som har extern politisk bärighet för bättre integrering och samordnad behandling av programmen .
Herr talman , herrar kommissionärer , kära kolleger !
Leader I var en verklig framgång , framför allt tack vare den flexibla administrativa förvaltningen mellan kommissionen och de lokala aktörerna .
Jag tycker att det är beklagligt att kommissionen inte upprättat samma bokslut över Leader II , ett bokslut över projektens kvalitet , mängden förbrukade anslag och framför allt över att vissa lokala aktörer givit upp inför den administrativa och ekonomiska tungroddhet man stött på .
Jag gläds emellertid åt att nya medel inrättats , inom ramen för Leader + , för att hjälpa landsbygdsområdena att utveckla sin potential och genomföra målsättningarna med lokal och hållbar utveckling .
Jag vill särskilt betona experiment med nya former för att förädla natur- och kulturarvet och förstärka den ekonomiska miljön , för att främja sysselsättningen .
Jag tror man kan anta att utbyte av dessa positiva erfarenheter av utvecklingen också kan förekomma inom ramen för det gränsöverskridande samarbetet .
Det är också intressant att notera att alla landsbygdsområden är stödberättigade enligt Leader II .
Om emellertid möjligheten kvarstår för medlemsstaterna att , inom ramen för detta initiativ , fastställa områden , bör kommissionen se till att det finns en viss koncentration av resurserna och prioritera projekt inom mindre framgångsrika områden .
Det krävs naturligtvis öppenhet om urvalskriterierna när det gäller projekt och lokala aktionsgrupper .
Det förefaller mig också som om man framför allt skulle behöva se till att staternas eller de lokala myndigheternas ekonomiska system inte längre är de som orsakar betalningsförseningar , något som försatt vissa lokala aktionsgrupper i konkurs inom ramen för Leader II .
Herr talman !
Som ledamot från ett yttre randområde måste jag säga att det är en mycket speciell eftermiddag när det gäller regionalpolitiken och det säger jag med anledning av debatten om två gemenskapsinitiativ , Urban och Interreg .
Jag vill påminna om att nämnda initiativ syftar till att , när det gäller det första , Urban , att förbättra livskvalitén för medborgare som bor i stadsdelar i olika europeiska städer , och Interreg , att främja sammanhållningen och att se regionernas mångfald och möjligheter i Europeiska unionen , särskilt när det gäller att inkludera de yttre randområdena i kapitel B och C. Vi beklagar , precis som föredraganden , att kapitel IIIA har tagits bort .
Vi anser att hänvisningen i Interreg att skapa ett europeiskt övervakningscentrum om samarbetets effekter är mycket klokt .
Tack till föredragandena , särskilt Decourrière för hans känslighet för de regionala frågorna och för att han accepterat våra ändringsförslag .
Jag hoppas att kommissionären godkänner det förslag vi lägger fram .
Herr talman !
När det gäller de olika initiativ vi behandlar denna eftermiddag vill jag strikt uppehålla mig kring en reflektion kring ett av dessa .
Det gäller rent konkret Urban-programmet .
Det är sant att vi i dag debatterar detta program eftersom Europaparlamentet envisades med att det skulle vara kvar .
Kommissionens förslag var att ta bort det , tillsammans med andra initiativ , men parlamentets förslag och kommissionens egen känslighet när det kom till kritan gjorde att Urban-programmet bibehålls .
Jag tycker att vi skall glädja oss över det .
Men , vilka var kommissionens argument , och i synnerhet kommissionär Monika Wulf-Mathies samt generaldirektör Eneko Landaburu , för att Urban-programmet inte skulle vara kvar ?
Argumentet var tungt .
Den urbana frågan är så viktig att vi inte kan begränsa den och nästan nedvärdera den med ett program som har en väldigt liten budget .
I dag har vi programmet och jag tror således att vi uppnått något viktigt , detta tecken på identitet som Urban är för Europeiska unionen .
Men jag skulle vilja vända mig till kommissionär Barnier för att lägga vikt vid kommissionärens och generaldirektörens argumentation eftersom jag tror att de hade väldigt rätt .
Den urbana dimensionen bör innefattas oerhört mycket djupare i alla strukturfonder .
Den budgetnivå våra städer behöver - där 80 procent av den europeiska befolkningen lever och som till stor del håller på att utvecklas till det goda och det dåliga vi har i Europa - , tror jag kräver att denna europeiska dimension beaktas och Urban-programmet får inte vara rättfärdigandet för att inte på djupet analysera , att inte prioritera och därför inte införa ett budgetanslag som vida överstiger det tidigare i program som påverkar städerna genom alla de europeiska fonderna .
Därför anser jag att det är onödigt att åter upprepa det antal faktorer som kräver denna investering i de urbana områdena , faktorer som är på dagordningen .
Jag skulle vilja förmedla till kommissionären att vi hoppas på förståelse för detta .
Samtidigt som vi välkomnar det sektorsövergripande förhållningssättet som finns i det nya Equal-initiativet , är det mycket viktigt att programmet behandlar de typiska former av diskriminering som i synnerhet skadar handikappade personer : Fysiska hinder på arbetsplatsen som påverkar dem med begränsad rörlighet , visuella informationssystem som inte är till nytta för blinda anställda , arbetssystem som effektivt hindrar dem som har inlärningsproblem eller psykiska problem .
Handikapporganisationer och handikappade personers icke-handikappade företrädare måste få lämplig insyn vid beslutsfattandets alla stadier .
Detta är skälet till varför detta parlament har lagt fram punkterna 10 och 15 i resolutionen för att se till att medlemsstaterna inte skall kunna bortse från någon målgrupp .
De handikappade har alltför ofta uteslutits från listan .
Eftersom handikappade inte utgör en enda homogen grupp - många döva ser t.ex. sig själva som en språklig minoritet som inte erhåller respekt för sitt eget språk och sin egen kultur - är det nödvändigt , vilket uttrycks i punkt 9 , att tillåta att vissa partnerskap bestäms som är specifika för ett särskilt handikapp eller en annan grupp .
Equal-initiativet är fortfarande mycket viktigt också i regioner som min hemregion i östra England , som i princip inte kan komma i fråga för stöd från mål 1-fonderna .
Vi har haft extra starka incitament för att erhålla medel från gemenskapsinitiativ och kan uppvisa en utmärkt historik .
Före detta Adapt-projekt som sträcker sig från Core-projektet - genom vilket man har utvecklat nya leverantörskedjor inom bilindustrin i Bedfordshire - till standardhöjande projekt för mindre företag i Hertfordshire i Essex .
Vi har sett hur Now-projektet har hjälpt 70 kvinnor att få arbete i Suffolk , av vilka många kunde komma och dela med sig av sina erfarenheter direkt med oss i Europaparlamentet i Bryssel .
Equal-initiativet är fortfarande viktigt för oss , eftersom det är just i relativt sett mer välmående regioner där icke-kvalificerade arbetstillfällen försvinner , och det är denna typ av arbeten som kan vara en viktig första hållplats för dem som är diskriminerade på arbetsmarknaden .
Till sist några ord om Interreg .
Egentligen är det rent nonsens att partnerskap som upprättats 1994 nu förlängs med undantag av nya interregionala förbindelser .
Under denna period har hamnarna Great Yarmouth och Harwich på Essex-Suffolk-Norfolkkusten infört betydelsefulla nya transport- och ekonomiska förbindelser med partner i Nederländerna .
Jag uppmanar parlamentet att stödja vårt ändringsförslag 2 , vilket kommer att säkerställa flexibilitet genom att inkludera nya områden , i synnerhet när det gäller havsgränser .
Herr talman , ärade kommission , ärade damer och herrar !
Herr talman , jag vill för allas information komma med ett klarläggande .
Förbundskansler Schüssels regering fortsätter driva förre förbundskansler Klimas socialdemokratiska regerings flyktingpolitik .
Det förekommer ingen ändring av flyktingpolitiken i Österrike !
Landsbygdsområdena utgör över 80 procent av EU : s yta , och 25 procent av befolkningen lever här .
Som bondkvinna och ledamot har jag alltid varit angelägen om att inte se jordbruket som något för sig , utan att se till hela landsbygdsområdet .
Särskilt värdesätter jag en integrerad satsning på landsbygdens utveckling eftersom jag är övertygad om att man kan skapa en aktiv och attraktiv livsyta för alla endast genom att sammanföra alla yrkesgrupper och alla människor på landsbygdsområdet till en gemenskap , kort och gott - landsbygdsområdets mångfaldiga funktion .
Det nya Leader + -programmet hälsar jag särskilt välkommet på grund av dess omfattande karaktär .
Det kommer i framtiden att bli möjligt att ha program inte bara i de enskilda stödområdena , utan i alla regioner inom EU .
Denna horisontella satsning är vettig i och med att programmen för landsbygdens utveckling också är utformade så .
Finansieringen kommer framdeles inte längre att skötas via tre fonder , utan då endast ur Europeiska utvecklings- och garantifonden för jordbruket ( EUGFJ ) .
Därför kommer det att krävas en höjning av kvalitén på programmen , för EUGFJ skall vara ett verksamt finansieringsinstrument .
Högre precision vid urvalet kommer att leda till höjd effektivitet , för pengarna skall inte slösas bort planlöst .
Jag vill också peka särskilt på den punkt som bildar en ansats till en integrerad och miljöanpassad utvecklingsstrategi .
Detta innebär att det finns en stor sysselsättningspotential för framtiden på landsbygdsområdet , och vi måste utnyttja detta om vi vill ge människorna på landsbygden ett perspektiv .
Därför är politik på landsbygden mer än politik bara för bönderna .
Leader + skall komplettera redan befintliga program , undvika överlappning och dubbelfinansiering och bidra till en så omfattande utveckling som möjligt .
På så sätt kan Leader + tillsammans med programmen i förordning 1257 / 99 backa upp andra stöttepelaren i den gemensamma jordbrukspolitiken ännu mer och åstadkomma bästa möjliga resultat för det samlade landsbygdsområdet .
Herr talman , bästa kolleger !
Jag är inte alltid stolt över vad det här parlamentet sysslar med , men Urban-programmet är ett av de bästa exemplen på vår verksamhet , det uppstod just på parlamentets initiativ .
Kommissionen ville avskaffa Urban , men den här gången drog parlamentet det längsta strået .
Det är bra att Urban fortsätter , ty man har på lokal nivå fått goda resultat av det .
Problemen i europeiska stadsområden håller på att bli värre ; som tur är delar vi nu åsikt med kommissionen .
Majoriteten av Europas befolkning bor i städer , deras problem är bland de viktigaste inom regionalpolitiken och mycket komplicerade frågor .
Risken för utslagning är stor .
I många franska och engelska städer finns redan slumområden där många onda ting föds .
Ingen av oss vill ha sydamerikanska favelas i Europa .
Vi måste agera nu innan det är för sent .
Städerna spelar också en avgörande roll för den europeiska ekonomin .
Vi återkommer alltid till samma europeiska grundproblem : vårt näringsliv är inte tillräckligt dynamiskt och uppmuntrar inte individen i tillräckligt hög grad .
Näringslivet måste vara starkt om vi skall kunna ta hand om våra närstående och vår miljö .
Detta är inte politik utan livets enkla logik .
När det gäller användningen av pengar är det bra att pengarna nu har centraliserats , ty om man sprider skotten åt alla håll försvinner krutet all världens väg som en flock sparvar .
Nu måste vi koncentrera oss på att lösa de små och medelstora städernas problem eftersom de inte har tillräckligt med kritisk massa .
På det sättet kan vi också ge mera fart åt de omgivande landsbygdsregionerna ; man glömmer ofta att städernas och landsbygdens problem i själva verket går hand i hand .
Grunden för allt är att man skall uppmuntra individens innovativa förmåga och företagsamhet eftersom den massrörelse som skapar en intern regional reform börjar hos en individ .
Att ge finansiering utan att det finns en ekonomi som står på egna ben är som att bära vatten till en sinad brunn : drickat räcker för en stund , men i morgon är brunnen åter tom .
Herr talman !
I och med att Interreg III förverkligas går den europeiska samarbetspolitiken in i en ny fas .
Vår uppmärksamhet riktas inte längre enbart mot de inre gränserna , utan även mot de yttre .
I dagens läge med globalisering och kulturell öppenhet behöver Europeiska unionen instrument för att stärka sina band och sina kommunikationskanaler med angränsande regioner , särskilt i Öst- och Sydeuropa .
Unionens gränser får inte längre utgöra ett hinder för en balanserad utveckling utan tvärtom en möjlighet , en bro till ett mer fruktbart samarbete .
Via de ändringsförslag som har antagits i utskottet försöker parlamentet komplettera kommissionens arbete genom att föra in nya namn på listan över mottagarområden för stöden , särskilt till förmån för de yttre havsgränserna i Sydeuropa .
I sitt förslag till riktlinjer påpekar kommissionen faktiskt att dessa gränser fordrar större uppmärksamhet än tidigare .
Detta med beaktande av utvidgningsprocessen mot öst och processen för större integrering med Medelhavsländerna .
Som ordförande Prodi också påminde om när han lade fram de strategiska målen för 2000-2005 är nylanseringen av Barcelonaprocessen en prioriterad fråga för unionen , och Interreg III-initiativet kan ge sitt bidrag till att detta strategiska mål uppnås .
Vi gläder oss åt det utmärkta arbete föredraganden har gjort och hoppas bara att kommissionen tar vederbörlig hänsyn till de förslag parlamentet har lagt fram , i enlighet med åtagandena i uppförandekoden för genomförande av strukturpolitik , och med de ändringar som behövs bekräftar detta gemenskapsinitiativs omvandling från att enbart vara ett instrument för intern omfördelning till att bli en möjlighet att nylansera och värdesätta relationerna med grannländerna .
Herr talman !
Från i år står runt 200 miljarder euro till förfogande för strukturfonden fram till år 2006 , men bara 5 3 / 4 procent har reserverats för gemenskapsinitiativen : Interreg , Leader , Urban och Equal .
Det är en minskning med 3 3 / 4 procent mot hittillsvarande gemenskapsinitiativ .
För Equal har inte mer än 2,8 miljarder euro avsatts , vilket framgår tydligt av kollegan Ursula Stenzels välbalanserade betänkande .
Desto mer förvånande är det stora antalet ändringsförslag och den långa önskelistan som rör möjliga uppgifter .
Hur skall man då prioritera ?
Det råder enighet om grundsatsen att diskriminering och ojämlikheter på arbetsmarknaden skall arbetas bort .
Transnationella strategier skall ge eftersatta grupper tillgång till sysselsättning .
Jag har ingen förståelse för förslag som innebär att man vill satsa på byråer för utbyte av information om tekniskt bistånd .
Dessa byråer var faktiskt föremål för den mest häftiga och berättigade kritik mot den förra kommissionens arbete .
Vårt utskott för sysselsättning och socialfrågor gick nu en gång i spetsen för analysen av väsentliga brister och försummelser i kontrollen av Leonardo .
Kommissionen kan således inte heller när det gäller Equal slippa undan det direkta ansvaret och kontrollen .
Förslag från medlemsstaterna kan kommissionen godkänna endast om dessa uppfyller alla villkor .
För det första : integreringsarbetet genom sektoriella och geografiska utvecklingspartnerskap , varvid hänsyn skall tas till sysselsättningspolitiska grundprinciper .
För det andra : systematisk integrering av berörda aktörer , de lokala , regionala och nationella myndigheterna , utbildningscentren , universiteten , de frivilliga organisationerna , arbetsmarknadens parter och den privata sektorn med ett bestående partnerskap som mål .
För det tredje : en garanterat entydigt innovativ karaktär på metoder och modeller .
Kommissionen måste alltså förpliktas vad gäller den strategiska ramen för att främja arbetsförmåga och arbetskvalitet , utvärdering av resultaten och den effektiva kommunikationen kring best practices .
Först då kan man uppnå den önskade multiplikatoreffekten .
Herr talman !
Jag vill hänvisa till kommissionens förslag om budgetposten för främjande av den gemensamma jordbrukspolitiken .
Den 26 oktober 1999 antog Europeiska kommissionen ett förslag för att se till att budgetposten för information till allmänheten om den gemensamma jordbrukspolitiken ( GJP ) får en rättslig grund .
Genom detta förslag kommer den befintliga budgetposten B2-5122 att tas bort och en ny budgetrubrik , B1-382 , kommer att skapas .
Åtgärder som främjar en förståelse mellan unga jordbrukare och EU , och som också skapar starkare förbindelser med ansökarländerna och resten av världen är viktiga .
Jag lägger därför fram dessa ändringsförslag i parlamentet för att detta skall ge sitt stöd till de bidrag som denna typ av program ger .
Med beaktande av behovet av att uppmuntra unga jordbrukare att fortsätta driva sin verksamhet , är det oerhört viktigt att de håller sig väl informerade om utvecklingen inom den gemensamma jordbrukspolitiken .
Information till och fortbildning av unga jordbrukare på gemenskapsnivå är oerhört viktigt .
Jag ber er att stödja att en del av den tillgängliga budgeten skall koncentreras på kunskapsutveckling bland gemenskapens unga jordbrukare .
Vad gäller information och fortbildning , så har denna budgetpost tidigare använts för tilldelning av medel till information , kommunikation och fortbildning .
Men kommissionen föreslår nu att fortbildning inte längre skall ingå .
Jag anser att fortbildning bör ingå i de fall denna ger relevant information om GJP på gemenskapsnivå .
En sådan fortbildning på gemenskapsnivå är ett sätt att se till att unga jordbrukare har den information om GJP som är nödvändig för att kunna fatta bra affärsbeslut för framtiden .
Jag lägger därför fram tre ändringsförslag .
Jag uppmanar parlamentet att stödja dessa .
Herr talman !
Jag tar till orda för att , med erfarenhet från den kommunala förvaltningen , uttrycka nyttan av , jag vågar säga nödvändigheten , att Urban-programmen har tre inriktningar .
För det första att främja återställande av historiska , gamla , kanske ödelagda infrastrukturer och stadsdelar .
För det andra att främja och stimulera den ekonomiska aktiviteten och det sociala livet i dessa historiska kvarter , i dessa delar av de gamla städerna .
Vi har ingen större nytta av gator , som nu kanske har utmärkt belysning , med nya trottoarer , med stenbeläggning , kanske vitkalkade och vackra , om vi inte har förmåga att fylla dem med aktivitet och således också sysselsättning .
Jag vill förtydliga att det inte handlar om finansiering eller hjälp till olika sociala aktörer utan att också finna en inriktning mot sysselsättning i urvalet av stödberättigade projekt eller , vilket är detsamma , projekt som leder till att gynna skapande av , impulser till och initiativ för sysselsättning .
För det tredje - och kanske skulle man behöva säga att det är det första - , att projektens huvudinriktning måste vara ett fullständigt återvinnande av personer och familjer , eftersom människan inte är gjord för rätten , utan rätten för människan .
I dessa områden i våra städer lever ofta ensamstående föräldrar , äldre som lever på pension och inte längre deltar i produktionen och familjer med svårigheter , ibland upplösta och ostrukturerade .
De bor i områden som borde kunna dra nytta av dessa projekt .
Om vi kan uppnå detta med dessa tre inriktningar tror jag att dessa familjer , dessa personer , dessa europeiska medborgare kommer att tro mer på Europa och det tycker jag är mycket viktigt eftersom det i slutänden är städerna som kommer att bli mer och mer huvudrollsinnehavarna i det europeiska samhällslivet .
Herr talman , herr kommissionär !
Det är i dag uppenbart att jordbruket i sig har allt svårare att behålla kvar befolkningen på landsbygden , speciellt ungdomar .
Den nyligen offentliggjorda sjätte periodiska rapporten om den sociala och ekonomiska situationen och utvecklingen i Europeiska unionens regioner pekar på just detta , och visar att de 25 jordbrukstätaste regionerna i Europeiska unionen är de som har högst arbetslöshetsnivå , förutom sina traditionella problem med en åldrande befolkning och utbredning av ödemark .
I detta sammanhang har kommissionen , undan för undan , tyvärr alltför långsamt , lagt fram initiativ som på sikt balanserar eller kompletterar den gemensamma jordbrukspolitiken , och strävar efter att omfatta en större del av landsbygdens resurser , och uppbåda dessa i initiativ och investeringar som gynnar befolkningens välfärd , oavsett de är jordbrukare eller ej .
Detta är fallet med den senaste utvecklingspolitiken för landsbygden som inleddes i Agenda 2000-reformen och det är särskilt fallet med gemenskapsinitiativet Leader som lades fram med Leader I och II , 1991 och 1994 , och som nu fortsätter i Leader + .
Jag skulle därför vilja understryka tre frågor : den första är att det är viktigt att urvalet av de lokala aktionsgrupperna ( GAL ) som ansvarar för organisationen och genomförandet av projekten , inte är politiska , och det bör ske ett urval enbart utifrån meriter för projektet och man bör prioritera dem som har arbetat mest i organisationer utanför myndigheterna , vilka i inget fall bör utgöra mer än 50 procent av partnerna i GAL ; den andra frågan är att i samarbetsåtgärderna mellan de lokala aktionsgrupperna och liknande organisationer i tredje land skall respektera kommissionens ursprungliga skrivning - punkt 18 - och inte den i Starkommitténs restriktiva version , som genomförts mot detta parlaments vilja .
Därför lade jag fram ett ändringsförslag i detta syfte , vilket utskottet för jordbruk och landsbygdens utveckling godkände och som jag hoppas kammaren godkänner ; för det tredje skulle jag vilja påminna om att det är nödvändigt att Leader , efter år 2006 , övergår från att bara vara ett gemenskapsinitiativ av pilotkaraktär till att också ta med utvecklingen av landsbygden i den gemensamma jordbrukspolitiken vilken enligt min åsikt borde byta namn till " den gemensamma jordbruks- , regional- och landsbygdspolitiken " .
Jag skulle vilja gratulera vår kollega Procacci till det utmärkta betänkande han har lagt fram . .
( FR ) Herr ordförande !
Innan mina kolleger och vänner , Franz Fischler och Anna Diamantopoulou , uttalar sig - eftersom vi haft turen att delta i denna debatt med samma uppmärksamhet alla vi tre som är ansvariga för dessa fyra gemenskapsinitiativ - , skulle jag vilja försöka ta upp Urban och Interreg , som många av er erinrat om .
Jag vill till att börja med framföra mitt tack till föredragandena från utskotten , från alla utskott , men också till gruppernas talare och till var och en av er för den stora kvalitet och det stora intresse som era inlägg vittnar om när det gäller dessa två initiativ .
Det gäller särskilt det som Arlene McCarthy sade om Urban , och jag vill tacka henne inte bara för det arbete och det betänkande hon lagt fram utan också , och varför skulle jag inte i min tur säga det , för det vi är skyldiga henne , för det ni är skyldiga henne när det gäller detta initiativ , liksom det vi mer eller mindre är skyldiga ert parlament .
Det är faktiskt Europaparlamentet som politiskt beslutat och önskat bibehålla detta initiativ , till förmån för förnyelse av städer som befinner sig i kris , till förmån för en hållbar stadsutveckling som samtidigt omfattar detta integrerade synsätt , som vi fäster stor betydelse vid , för att behandla såväl ekonomiska som sociala och miljömässiga aspekter .
Andra punkter där vi är överens , och som betonats i Arlene McCarthys betänkande , är hur effektivt detta instrument är , tack vare den ekonomiska koncentrationen och den kritiska nivån för ingripandena , den horisontella mekanismen , som tycks vara gynnsammare för att sprida resultaten och öka utbytet av erfarenheter och goda tillämpningar , och slutligen de lokala myndigheternas ökade betydelse när det gäller utformning och förvaltning av programmen , på grundval av ett verkligt partnerskap .
Efter att ha erinrat om de grundläggande punkter där kommissionens och parlamentets förslag är samstämmiga och efter att ha betonat att jag tyckte det var mycket intressant att lyssna till de olika inläggen , skulle jag nu vilja besvara viss kritik , mot vissa förslag som lämnats , och jag ber om ursäkt i förväg för att jag inte kan citera varje talare personligen .
Jag tror emellertid att de kommer att känna igen sig .
Programmet Urban , till att börja med , och maxtröskeln med femtio städer , som vissa av er bedömt som godtycklig .
Jag förstår denna oro .
Jag har därför bett mina enheter att överväga en rimlig ökning av antalet städer som kan vara berättigade till stöd från Urban , med hjälp av vissa garantier om koncentration , till att börja med - jag tänker bl a på områden för åtgärder som måste omfatta minst 20 000 invånare och undantagsvis 10 000 invånare - och sedan också på den kritiska ekonomiska massan : vi måste hålla oss till 500 euro per invånare för att Europeiska unionens åtgärd skall vara både effektiv och begriplig , och för att den inte skall likna någon fördelning av anslag mellan flera mottagare , som inte längre skulle vara begriplig för medborgarna eller kommunerna .
Det var mitt första svar på frågan om tröskeln .
När det gäller den andra frågan , som handlar om kompletterande kriterier som borde beaktas vid urval av områden med svårigheter , är jag också här beredd att visa prov på större flexibilitet och överväga andra relevanta kriterier , som komplement till gemenskapens kriterier i punkt 11 i förslaget till riktlinjer .
Punkt tre : särskilda åtgärder till förmån för vissa socialgrupper - flera av talarna har erinrat om detta - kvinnorna , men också invandrarna , flyktingarna , borde tas med .
Mina damer och herrar parlamentsledamöter !
Denna oro står i centrum för vårt initiativ Urban och om det är nödvändigt är jag beredd att eventuellt skriva om texten så att budskapet skall bli ännu tydligare .
Jag skulle när det gäller Urban vilja avsluta med att tala om villkoren för genomförande , och till att börja med urvalsförfarandet .
Vissa har önskat att det skulle vara mindre byråkratiskt , mer öppet , att vi skulle undvika onödig användning när det gäller projekt och finansiering .
Mina damer och herrar !
På denna punkt måste vi vara tydliga : enligt subsidiariteten är urvalet av stödberättigade områden eller kommuner för Urban framför allt medlemsstaternas ansvar .
Kommissionen är för sin del beredd att undvika all omotiverad byråkratisk överbelastning , men vi kan inte - och ni kanske skulle vara bland de första att förebrå oss det - avstå från att kontrollera relevansen och kvaliteten i de program som föreslås .
Den andra anmärkningen gäller tidsfristen för att lämna in program , och möjligheten att lägga fram kompletteringar till programplaneringen tillsammans med programmen .
Jag har inga invändningar mot denna idé om att överlämna ett komplement till planeringen tillsammans med huvudprogrammet .
Detta får emellertid inte innebära att den ursprungliga tidsfristen förlängs .
Jag erinrar om att den är sex månader för detta program .
Denna tidsram , som för övrigt är identisk med den som vi beviljat för Interreg och för samlade programplaneringsdokument inom mål 2 , borde i allmänhet vara tillräcklig för att upprätta ett program , tycker jag , vilket inte hindrar att projekten definieras senare .
När det gäller Urban skulle jag vilja avsluta med en sista kommentar .
Någon av er önskade att denna stadsdimension inte bara skulle begränsas till Urban .
Det instämmer jag helt i .
Jag berättade själv vid mötet med ministrarna för fysisk planering och stadsplanering om min oro - och jag är verkligen oroad - över att stadsaspekten i samlade programplaneringsdokument och gemenskapsstödramar , i de programplaneringar där vi inleder förhandlingar , skall hamna utanför Urban , bland alla program inom mål 1 och mål 2 , och jag tror att jag kan påstå att vi är vaksamma , men att man också kan utläsa denna stadsdimension utanför Urban i hela programplaneringen av strukturfonderna .
Men för framtiden , för vi måste ju se framåt , är jag mycket angelägen om att se hur Urban konkret kommer att genomföras , och jag är också mycket angelägen att se vilken erfarenhet eller vilka lärdomar vi kan dra , eftersom denna stadsdimension uppenbarligen kommer att stå i centrum för vad som , i den kommande budgetplanen , skulle kunna vara en ny europeisk politik för fysisk planering .
Jag glömmer inte , vi kan inte glömma , att 80 procent av de europeiska medborgarna i dag lever i städer och det är anledningen till att Urban är mycket viktigt .
Jag upprepar på nytt att vi måste vara uppmärksamma på stadsdimensionen i hela programplaneringen för strukturfonderna .
Herr ordförande !
Jag skulle nu vilja ta upp Interreg och , precis som jag gjorde när det gällde Arlene McCarthy , tacka er föredragande , Francis Decourrière , för ett bra och relevant arbete .
Han har betonat flera punkter där både vi och flera av er kan instämma : betydelsen av detta transeuropeiska samarbete , med dess tre områden , gränsöverskridande , transnationellt och interregionalt , det mervärde som Interreg medför för gemenskapen , hur begripligt det är jämfört med den allmänna ramen för strukturfonderna , och den verkligt gränsöverskridande och transnationella förstärkningen av programmen och de stödberättigade åtgärderna , betydelsen av gemensamma strukturer - det som jag , apropå en annan debatt som börjar i dag , nämligen regeringskonferensen , kallat européernas gemensamma anda som vi måste förstärka , med Interreg och tack vare Interreg , hur vi skall förstärka den gemensamma andan via gemensamma strukturer för genomförande av programmen med verklig ekonomisk solidaritet , betydelsen av partnerskapet för att garantera aktivt deltagande i alla berörda lokala och regionala myndigheter samt föreningar inom den privata sektorn och sociala och ekonomiska partnerskap .
Efter dessa allmänna kommentarer skulle jag vilja koncentrera mitt inlägg beträffande Interreg på era huvudsakliga kommentarer .
De första gäller tidsfristen och innehållet i detta initiativ .
Ni säger att antagandet av dessa riktlinjer skett alltför sent , och risken att tidigare program skulle avbrytas har betonats , bl.a. av er föredragande .
Det är sant , det erkänner jag , och ni vet mycket väl orsakerna , mina damer och herrar parlamentsledamöter .
Antagandet av riktlinjerna för Interreg är försenat till i mars-april 2000 .
Jag erkänner det , jag noterar det precis som ni .
Jag noterar emellertid också att medlemsstaterna och regionerna redan aktivt förbereder programmen för Interreg III , och förslaget till riktlinjer har för övrigt redan delats ut för mer än tre månader sedan .
Jag noterar också att utgifterna blir stödberättigade så snart programmen lagts fram och jag bekräftar att principen med retroaktivitet kommer att gälla ända till den 1 januari , om programmet läggs fram före den 30 april .
Så långt min första kommentar .
Kommentar två : när det gäller den ofullständiga förteckningen över åtgärder inom område B vill jag bekräfta att jag bett kommissionen att acceptera att andra specifika teman införlivas , bl.a. till förmån för små och medelstora företag eller kulturarvet , i förteckningen över åtgärder som kan vara stödberättigade inom område B , och att man alltså inte skall betrakta denna förteckning som fullständig .
Punkt tre gäller samarbetet mellan regioner , och betydelsen av område C. Kommissionen instämmer i kammarens kommentarer om betydelsen av område C för samarbete mellan regioner .
Enligt er föredragandes önskemål skall jag överlämna detaljerad information till er om systemet för att genomföra detta område .
Kommentar fyra gäller övervakningscentrum och eventuellt utnyttjande av ett kontor för tekniskt bistånd .
Såsom ni begärt har jag beslutat att ta bort alla hänvisningar till ett kontor för tekniskt bistånd i texten , i avvaktan på att den pågående debatten inom kommissionen om systemen för att utlokalisera enheterna får en lösning .
Mina damer och herrar parlamentsledamöter !
Om vi avskaffar alla hänvisningar till och senare allt utnyttjande av ett kontor för tekniskt bistånd får det konsekvenser , nämligen att antalet tjänster måste utökas för att utföra detta arbete , eftersom någon ju måste göra det , och man inte i evighet kan omstrukturera samma personal , även om våra uppgifter ökar med Ispa och med strävan efter att med större stramhet och öppenhet kontrollera gemenskapens anslag , som jag är ansvarig för , ofta i partnerskap med medlemsstaterna eller med dem som medansvariga .
När det sedan gäller genomförandet av Interreg , ett ämne som tagits upp av flera av er , och det eventuella stödberättigandet under område A , " gränsöverskridande samarbete " , åtgärder i Adriatiska havet , för Sicilien eller de yttersta randområdena , förstår kommissionen er oro och uppfattar tydligt er begäran under dessa olika punkter , mina damer och herrar .
Jag har därför för avsikt att ändra riktlinjerna för att i det gränsöverskridande området B införliva en specifik prioritering : " Integrerat samarbete för havs- och öregionerna " , för att vi på ett lämpligt sätt skall kunna täcka de olika möjligheterna till samarbete mellan dessa regioner .
Detta är en första öppning tillsammans med andra som vi redan föreslagit medlemsstaterna : större ekonomisk flexibilitet mellan område A och område B. Tack vare dessa två öppningar kan jag säga att kommissionen är beredd att granska fallet med de italienska regionerna och regionerna i tredje land vid Adriatiska havet , för att främja det mest lämpade samarbetet inom ramen för Interreg , och även med andra instrument , så snart dessa blir tillgängliga .
Jag har avslutningsvis beslutat att de yttersta randområdena , som jag är särskilt mån om , särskilt prioriteras inom ramen för det gränsöverskridande området i Interreg , med en samarbetsstrategi för att förbättra förbindelserna med deras grannländer och andra regioner i medlemsstaterna .
Jag vill också säga att jag är mycket mån om ett gott samarbete mellan Interreg och Europeiska utvecklingsfonden , bl.a. när det gäller Västindien och Indiska oceanen .
Allt detta borde göra det möjligt för oss att , utöver anslagen inom mål 1 och tillsammans med dem , bekräfta unionens roll som " aktiv gräns " .
Jag instämmer i den politiska målsättningen att unionens sju yttersta randområden verkligen skall vara unionens aktiva gränser , även om och just för att de ligger långt bort och är belägna i andra regioner i världen , där vi bör ha inflytande och vara aktiva .
En annan punkt jag vill ta upp är samordningen mellan Interreg , Phare , Tacis och Meda .
Det stämmer att också där , och det erkänner jag objektivt , kvarstår verkliga juridiska svårigheter .
Jag vill inte förringa dem , men framsteg pågår för samarbete inom område A med kandidatländerna , även om svårigheterna i anslutning till förvaltningsförfarandet och till projektens omfattning kvarstår .
Kommissionen måste fortsätta på den vägen .
Jag skall personligen se till det .
En första gemensam kommitté för Phare / gemenskapsinitiativ kommer att äga rum under februari för att gå igenom denna samordning , och jag vill bekräfta för er att jag tillsammans med mina kolleger Verheugen , Patten och Poul Nielson är vaksam och tillgänglig i det hänseendet .
När det gäller tekniskt bistånd , avslutningsvis , där er föredragande och flera av er haft kommentarer , är det självklart att kommissionen skall följa bestämmelserna i artikel 23 i den allmänna förordningen om tekniskt bistånd , om det verkligen handlar om bistånd som utformas som ett instrument som kan användas för strukturpolitiken i allmänhet .
Enligt den allmänna förordningen skall emellertid alla åtgärder för tekniskt bistånd , som kan åberopa en viss koppling till ett gemenskapsinitiativ , föreslås enligt artikel 20 , och inte artikel 23 .
Det innebär att taket på 0,25 procent enligt artikel 23 inte är tillämpligt när det gäller detta slag av bistånd .
Mina damer och herrar !
Jag sätter stort värde på att vi , i vår strävan efter stramhet och öppenhet , ändå behåller vissa ekonomiska områden för allt som gäller utbyte av erfarenheter och information , men inte propaganda , och för att inrätta nätverk som garanterar god kommunikation mellan de bästa tillämpningarna inom unionen .
Min slutsats om Interreg , herr talman , mina damer och herrar , är att dessa gemenskapsinitiativ , som jag är ansvarig för , motsvarar ett verkligt behov och det som sagts här visar det .
De förebådar också en verklig europeisk politik för fysisk planering inom vår utvidgade union .
Kommissionen sätter därför , precis som ni , stort värde på detta .
Jag står till ert förfogande för att överlämna den tidigare översikten över programplaneringen som ni bett om , men också för att regelbundet hålla er informerade om genomförandet av dessa initiativ under den nya programplaneringsperioden .
Jag tackar återigen var och en av er , och särskilt Arlene McCarthy och Francis Decourrière , och jag skulle när det gäller dessa två initiativ vilja säga att de ligger inom en ekonomisk ram som ni känner till väl : bara 700 miljoner euro för Urban , men det är ändå bättre än ingenting , 4 miljarder 800 miljoner euro för Interreg .
Vi arbetar alltså inom denna ram och inte utanför den .
När det därför gäller dessa två initiativ vill jag , för att förtydliga de framtida strategiska och politiska diskussionerna inom fysisk planering och den kommande budgetplanen , framhäva att vi funnit denna konstruktiva dialog med parlamentet och dess utskott mycket intressant .
Det jag nu kunnat säga , mina damer och herrar parlamentsledamöter , visar att kommissionen är fast besluten att ta hänsyn till detta .
( Applåder ) Fru talman , ärade ledamöter , mina damer och herrar !
Låt mig inleda med att rikta mitt tack till herr Procacci för det betänkande som han har utarbetat .
Men jag vill också tacka alla berörda utskott och parlamentet för det breda stöd som man har gett initiativet Leader + .
Initiativet syftar till att ge landsbygdsområdet nya impulser att utveckla och utprova nya och originella satsningar , satsningar som sedan skall föras in som modell i allmänna program .
Jag är också glad att parlamentet i allt väsentligt stöder kommissionens uppfattning om att Leader + skall tillämpas i alla landsbygdsregioner , att överordnade prioriteringar skall införas och framför allt att även det aktiva samarbetet och sammanlänkningen mellan de olika landsbygdsområdena skall främjas .
Jag kan därtill konstatera att parlamentet delar kommissionens uppfattning att tillämpningen av Leader + följaktligen skall prioriteras i form av globala bidrag .
För att gå in på vissa detaljfrågor som har kommit upp här kan jag även bekräfta att vi vill ha så långtgående partnerskap och deltagande som möjligt för Leader + .
De olika grupperna , det må vara miljöorganisationer eller grupper som arbetar för sysselsättning , har möjlighet att medverka när kommissionen drar upp riktlinjerna .
Och det kommer inte heller att bli mindre , utan mer kapital som ställs till förfogande än under innevarande period .
Jag vill också påminna om att det inte är något nytt att vi inrättar ett övervakningscentrum .
Detta övervakningscentrum fanns redan för Leader I och Leader II .
Centrumet syftar uteslutande till att hålla igång just sammanlänkningen av de enskilda Leader-grupperna .
Finansieringen av övervakningsscentrumet får inte överstiga 2 procent av Leader-anslagen .
Vad gäller möjligheterna för projekt som har träning och utbildning som innehåll vill jag påpeka att just detta är en punkt som vi nu har integrerat i den nya utvecklingspolitiken för landsbygden , varför det i våra ögon inte längre är nödvändigt att göra så inom ramen för Leader .
Nu till innehållet i själva betänkandet .
Under punkt 14 uppmanar parlamentet kommissionen att omgående komma med en rapport om utvärderingen av Leader II .
Jag vill bara göra er uppmärksamma på att detta inte är särskilt meningsfyllt i nuläget eftersom kapital från Leader II ju fortfarande - och det ända till utgången av år 2001 - kan komma att redovisas .
Därför anser vi att det vore vettigare att genomföra denna utvärdering först när programmet har avslutats .
Naturligtvis kommer vi att göra detta och även se till att en rapport kommer er till handa .
Under punkt 18 föreslår parlamentet att ett kompendium över exempel på lyckade initiativ skall ges ut .
Jag kan bara tillägga att ett sådant redan finns .
Det har utarbetats av kommissionen och jag ställer det gärna till förfogande för alla intresserade ledamöter i kammaren .
Under punkt 21 betonar parlamentet att godkännandet av direktiven till Leader + från och med nu måste skyndas på för att programmen skall kunna köras igång .
Denna begäran stöder jag fullt ut .
Så snart yttrandet har godkänts här i parlamentet kommer riktlinjerna för Leader + ånyo att läggas fram i star-utskottet så att medlemsstaterna kan bekräfta det preliminära godkännande som man gav den 14 november .
Jag utgår från att kommissionen sedan kommer att kunna anta den slutgiltiga versionen av riktlinjerna i mars / april .
Och så snart dessa har offentliggjorts i Europeiska gemenskapernas officiella tidning återstår endast månaderna , nämligen de sex månaderna , för inlämning av förslag till Leader + -program .
Jag tycker det är viktigt att betona en sak : stöd kan utbetalas för Leader + från och med det datum då programmet kommer kommissionen till handa .
För de program som lämnas in före 30 april i år finns möjlighet att fastställa startpunkten för bidragsperioden retroaktivt till den 1 januari .
Under punkt 20 slutligen innehåller förslaget till resolution sju konkreta ändringsförslag för riktlinjerna .
Efter ingående prövning kan jag meddela att förslagen under punkterna 2 , 4 , 5 och 7 är godtagbara för kommissionen och kommer att antas .
Likaledes kommer förslaget under punkt 6 delvis att godkännas eftersom det bekräftas att fristen för att bevilja programmen inom Leader + uppgår till högst fem månader .
Ändringsförslaget under punkt 1 har i våra ögon hunnit bli inaktuellt i och med att punkten redan har omformulerats i parlamentets anda i anslutning till samrådet med representanterna för medlemsländerna i ansvariga utskott .
Följaktligen återstår endast ändringsförslaget under punkt 3 .
Kommissionen kan bara ansluta sig till denna begäran om ändring , för det överensstämmer exakt med kommissionens ursprungliga förslag .
Jag måste dock tillägga att våra aktionsgruppers samarbete med likvärdiga grupper i tredje land har gått för långt för medlemsstaterna .
Därför har vi fått en ändring i utskottet , men kommissionen kommer nu i den omarbetade versionen att ta hänsyn till parlamentets begäran på nytt och utforma riktlinjerna i enlighet därmed .
Kommissionen kommer även att kämpa vidare för att detta skall kunna godtas av medlemsstaterna .
I korthet om de 13 ändringsförslag som har lagts fram .
Här är det endast tre förslag som kommissionen inte kan godkänna , nämligen ändringsförslagen 3 , 12 och 13 .
Alla övriga kan kommissionen godkänna antingen fullt ut eller efter andemeningen .
( Applåder ) .
( EL ) Fru talman !
Damer och herrar ledamöter !
Det är ett egendomligt sammanträffande att vi i dag diskuterar Equal-initiativet här i Europaparlamentet .
I Europa har det den senaste tiden , på grund av den politiska utvecklingen i Österrike , funnits en stigande , en ökande politisk oro , det har gjorts politiska uttalanden och förekommit politiskt samtal .
Det bör betonas att såväl parlamentet som kommissionen har lagt fram särskilda strategier .
Särskilda förslag såväl om lagstiftning som om åtgärdsprogram som avser bekämpningen av diskriminering , som avser uppbyggnaden av samhällen med friheter och lagar .
Så , jag nämner helt kort paketet mot diskriminering och ber med anledning av det att de respektive ansvariga parlamentsutskotten utser föredragandena , så att vi så snabbt som möjligt kan gå vidare med paketet mot diskriminering .
Och jag kommer till Equal-initiativet , som naturligtvis grundar sig på artikel 13 .
Equal-initiativet avser alla former av diskriminering på grundval av artikel 13 , det vill säga bekämpning av diskriminering som grundar sig på ras , kön , ålder , handikapp .
Jag skulle särskilt vilja tacka Stenzel , för hennes arbete med att försöka nå en överenskommelse om Equal-initiativet är enastående svårt och komplicerat , såväl på grund av att utskott som ser på saken ur en annan synvinkel är inblandade som på grund av att det är en enastående känslig politisk fråga .
Min första kommentar , som även har formulerats av många kolleger , gäller frågan om huruvida kvinnorna måste tas upp separat .
Jag håller med om att det i artikel 13 finns en sak som vi inte håller med om , men fördraget är sådant i dag , och bland diskrimineringskategorierna finns på lika bas även diskriminering som grundar sig på kön .
Med fördraget som grund , i den form som det har i dag , är Equal-initiativet sammansatt på det sättet .
Jag vill dock påminna om att det finns en särskild pelare i sysselsättningsstrategin som gäller kvinnorna och att ett särskilt program , det femte programmet för jämlikhet mellan män och kvinnor , håller på att förberedas .
Jag har indelat frågorna som damerna och herrarna parlamentskolleger har berört i fyra grupper För det första , utvidgningen av de tematiska enheterna .
Det finns fyra tematiska enheter , liksom i sysselsättningsstrategin : anställbarhet , företagaranda , anpassningsförmåga och lika möjligheter , och vi instämmer i utvidgningen av dessa tematiska enheter i enlighet med de förslag som har lagts fram av Europaparlamentet .
Angående oron över risken att ett land lägger alla pengar på en av de kategorier som är utsatt för diskriminering , skall jag säga att det klart och tydligt sägs i initiativet att medlemsstaterna bör presentera en tematisk kategori för var och en av de grupper som är utsatta för diskriminering .
Den andra frågan gäller flexibilitet och förenkling .
Jag håller med Leinen om att språket i initiativet verkligen är mycket svårt och ogenomträngligt .
Av den anledningen håller avdelningarna redan nu på att revidera texten , att förenkla dess struktur och göra dess språk mer lättförståeligt .
Angående frågan om flexibilitet , vill vi med vårt förslag få till stånd utvecklingspartnerskap och utvecklingssamarbete , såväl på geografisk nivå , där grupper av olika slag skall samarbeta i en bestämd geografisk region för att bemöta diskriminering på arbetsområdet , som på tematisk nivå , där det till exempel skall kunna förekomma samarbete i en konkret ekonomisk sektor .
Här kommer det att finnas ett stort utrymme för flexibilitet i medlemsstaterna , och de kommer att kunna anpassa utvecklingssamarbetet i enlighet med sina önskemål .
En förutsättning är naturligtvis att medlemsstaterna samarbetar och att vi har ett nät med vars hjälp vi kan utbyta erfarenheter .
Avslutningsvis skall jag ta upp det tekniska biståndet .
Vi vill att det skall finnas fyra stödkategorier .
För det första skall förberedelserna stödjas , för det andra genomförandet , för det tredje samarbetet mellan aktörerna , så att ett erfarenhetsutbyte kommer till stånd , och för det fjärde det tekniska biståndet .
Eftersom det har funnits ett stort engagemang och en stor oro över frågan om hur det tekniska biståndet skall tillhandahållas , skall vi säga att externa byråer kommer att användas .
Det är omöjligt , vilket också min kollega Barnier sade , att kommissionens tjänstemän skall utföra allt det arbete som fram till i dag har utförts av externa medarbetare .
Målet är att det på nationell och europeisk nivå skall finnas stora grupper av åtgärder som offentliggörs , och det kommer att finnas en fullständig beskrivning av det arbete för vilket det externa biståndet begärs och en fullständig beskrivning av den produkt som vi förväntar oss av varje teknisk byrå , så att det är möjligt att både övervaka och utvärdera detta arbete .
Jag vill understryka att det är enastående viktigt att det aktuella initiativet främjas så snabbt som möjligt , dels på grund av politiska omständigheter , men även på grund av att vi anser att det är viktigt att det träder i kraft som planerat , dvs. att vi måste vara helt förberedda i slutet av 2000 .
Tack , fru kommissionär .
Jag skall till mina kolleger inom presidiet och berörda utskott framföra att ni gärna vill ha en snabb nominering av föredragande för de ärenden ni nämnde .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
( Sammanträdet avslutades kl .
20.40 . )
