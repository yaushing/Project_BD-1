 
Justering av protokollet från föregående sammanträde Protokollet från i går har delats ut .
Finns det några synpunkter ?
Herr talman !
Det står att jag röstade " för " Cunhas betänkande om fiske , när min avsikt var att rösta " emot " .
Jag vill gärna att protokollet rättas .
Och i debatten om Kina i går röstade jag för betänkandet .
Jag vill gärna att det tas med i protokollet .
Detta skall tas med i vederbörlig ordning , Wyn .
Herr talman !
Jag vill bara framkasta en fråga .
I gårdagens protokoll står det att vi diskuterat McNallys betänkande och att omröstning sker den 2 februari .
Jag vill bara fråga varför det måste vara så .
Jag har hört att det är något som inte stämmer med dokumenten .
Något sådant borde dock egentligen inte få ske .
Betänkandet har diskuterats , och vi hade i dag hunnit rösta om det , och jag förstår absolut inte varför en omröstning måste göras så långt efter debatten .
Kammarens princip har i sig varit att omröstningen bör genomföras så snart som möjligt efter debatten .
Anledningen till att vi skall genomföra omröstningen i februari är att vi har problem med vissa översättningar och detta måste vi lösa .
Vi måste ha överensstämmelse mellan de olika texterna och detta tar litet tid .
Det är ett rent tekniskt problem som uppstått på grund av översättningarna .
Herr talman !
Jag tog upp en sak i protokollet redan i går kväll .
Under punkt 6 i protokollet , på sidorna 6-7 , nämns mitt förslag om att punkt 6 i Cunhabetänkandet inte kan godtas .
Jag begärde en omröstning med namnupprop och talmannen förklarade tydligt att det skulle bli en omröstning med namnupprop om det .
Vi röstade också med hjälp av våra omröstningsmaskiner .
Men vad jag förstår har omröstningen inte registrerats .
Jag vill att det skall noteras att en omröstning med namnupprop borde ha ägt rum och att det borde ha funnits en förteckning med namnen på de som röstade för och emot förslaget .
Herr MacCormick , ordförandeskapet är medveten om det här problemet .
Det begicks dock ett ofrivilligt misstag , det vill säga den ansvariga personalen gjorde ett misstag som var absolut oförutsett , ofrivilligt , oundvikligt och helt omöjligt att förutse .
Så trots att omröstningen med namnupprop genomfördes korrekt så registrerades inte resultatet .
Det finns ingen annan anledning och det finns ingen möjlighet att lösa problemet .
Det är ödets nyck , MacCormick .
Herr talman !
I samma punkt , punkt 6 i gårdagens protokoll om förslag som rör förfaranden om Cunhabetänkandet , står det att jag återförvisade ärendet till utskottet enligt punkt 144 i arbetsordningen , främst för att det rådde tvivel om huruvida punkt 6 var tillåtlig .
Detta är inte korrekt .
Även om jag nämnde möjligheten av att min kollega MacCormick kunde väcka förslag om otillåtlighet , var skälet för en återförvisning till utskottet att det fanns betydande politiska motsättningar och praktiska oklarheter kring förslaget .
Jag ville därför ha ytterligare diskussioner och överläggningar med berörda parter .
Er anmärkning är noterad herr Hudghton .
Herr talman !
Jag har inga problem med vad som står i protokollet - det är vad som inte står i protokollet som är ett problem för mig .
I onsdagens protokoll finns en förteckning över ledamöter som har ändrat sin röstning .
Jag ser att det i gårdagens protokoll inte finns någon sådan förteckning , trots att jag känner till minst två ledamöter som ändrade sin röstning om resolutionen om kapitalskatt .
Jag vill gärna veta när vi får besked om dessa röstningsändringar , eftersom detta självklart är av intresse för vissa ledamöter .
Jag antar att ett tillägg kommer att göras till nästa protokollomgång , och att vi då får tillfälle att yttra oss .
Herr Ford , vi skall titta på detta och stämmer det så skall protokollet rättas i vederbörlig ordning .
Herr talman !
Jag vill bara informera er om följande : I morse förövades ett attentat i Madrid .
En bomb hade installerats i en bil .
En person har dött .
Jag vill bara å min grupps vägnar än en gång fördöma dessa terroristhandlingar .
Tack så mycket , fru Fraga .
Vi har faktiskt blivit informerade om den tragiska händelsen .
Än en gång bestraffas tyvärr det spanska samhället av dessa mordiska terrorister .
Ordförandeskapet noterar era ord med särskild intensitet eftersom ordförandeskapet vid dagens sammanträde också är spanskt .
( Protokollet justerades . )
 
Den gemensamma fiskeripolitiken : förstärkt dialog med industrin och andra berörda Nästa punkt på föredragningslistan är debatten om betänkande ( A5-0094 ) av Miguélez Ramos för fiskeriutskottet om förslaget till rådets förordning om förstärkt dialog med industrin och dem som berörs av den gemensamma fiskeripolitiken ( KOM ( 1999 ) 0382 - C5-0145 / 99 - 1999 / 0163 ( CNS ) ) . .
( ES ) Herr talman !
Med den förordning vi i dag granskar försöker man förstärka dialogen med industrin och andra berörda för den gemensamma fiskeripolitiken .
Kommissionen vill därmed försäkra sig om att informationen om yrkessektorns behov verkligen når fram och samtidigt underlätta en spridning av normgivande regler och gemenskapsbeslut inom ramen för fiskeripolitiken .
Fiskeriutskottet stöder givetvis det här förslaget till förordning .
För att kunna utforma förslag och utöva sina befogenheter behöver Europeiska kommissionen få lära känna verkligheten genom en dialog med de yrkesmän som ingår i denna .
Förslaget till förordning föregicks av en reform av den rådgivande kommittén för fiske och jordbruk , ett rådgivande organ som inrättades 1971 , och där alla yrkesgrupper ingår .
Sammanfattningsvis innebar reformen att nämnda organ aktualiserades genom att man införlivade andra huvudaktörer som under senare år har kommit att spela än allt viktigare roll i hanteringen av en förnuftig utvinning av resurserna , som till exempel de icke-statliga organisationer som är aktiva inom olika utvecklingsområden , miljöföreningar , konsumenter samt vetenskapsmän .
Reformen förde också med sig att sektorer som förut var underrepresenterade fick en större plats - fiskeodlingen samt marknadsföringen av produkterna .
Man ändrade även på antalet kommittéledamöter i plenum och specialiserade arbetsgrupper inrättades .
Jag skulle vilja säga att kärnpunkten i reformen av den rådgivande kommittén är att man nu prioriterar de organisationer som är representerade på gemenskapsnivå , så att kommittén inte bara blir ett språkrör för nationella ståndpunkter .
Parlamentets fiskeriutskott , och framför allt jag som föredragande för betänkandet , har starkt kritiserat det faktum att kommissionen inte rådfrågade oss när kommittén reformerades .
Detta innebär att vi i dag måste begränsa oss till att avge ett yttrande om förslaget till förordning , enligt min mening för litet .
När det gäller de mera konkreta områdena i kommissionens förslag att främja spridandet av information om den gemensamma fiskeripolitiken , de mål , mekanismer och lagbestämmelser som berör sektorn , så stöder vi dem till fullo .
Beslutar sig kommissionen för att driva igenom dessa informativa bemödanden så skulle inget , ärade kollegor , göra oss gladare .
Vid kommissionärens sista inställelse inför kommissionen erkände han att det var absolut nödvändigt .
Fischler sade att vi har problem med marketing och att det är nödvändigt att informera och värna om vår modell .
Intern information - mot den egna sektorn , inom vilken man ofta inte känner till eller är felinformerad om sin egen verklighet - samt extern information .
Som ledamot i fiskeriutskottet har jag många gånger förvånat mig över den stora okunskap som allmänheten har när det gäller den gemensamma fiskeripolitiken som är av stor vikt för många medlemsländer och för unionen i sin helhet .
När det gäller den interna informationen , till den egna sektorn , uppmanar vi kommissionen att ta hänsyn till den verklighet som många fiskare lever i .
Ärade kollegor , inte alla har tillgång till den nya tekniken och därför måste informationen och kampanjerna använda sig av alla medel som står till buds , inklusive de mer traditionella .
Här vill jag uppmärksamma tidskrifternas arbete - som oroar sig alltmer för det framtida fisket i Europa - liksom radio och TV , demokratiska instrument inom räckhåll för alla .
Avslutningsvis vill jag uppmärksamma kommissionen på representativiteten i de organisationer som ingår i den rådgivande kommittén .
Dialogen mellan kommissionen och yrkesmännen är väsentlig .
För att dialogen skall bli givande måste dock de yrkesmän man samtalar med verkligen företräda de olika sektorerna i den gemensamma fiskeripolitiken .
Varken i kommissionens förslag eller i regleringen av den rådgivande kommittén har man dock förutsett att det är så det skall vara .
I en så pulveriserad sektor , med enorm geografisk spridning men liten medlemsanslutning , riskerar man att kommissionens samtalspartner på gemenskapsnivå inte företräder de olika sektorerna på ett trovärdigt sätt .
För att öka representativiteten och komplettera vidtagna åtgärder så vore det kanske bra om kommissionen tog vissa initiativ för att stimulera en anslutning till de branschorganisationer som för närvarande finns .
Sektorns företrädare , som utsetts till kommissionens samtalspartner , med andra ord ledamöterna , är tvungna att företräda det gemensamma intresset .
Herr talman !
Jag stöder i stor utsträckning vad Miguélez just så modigt har framfört .
Ty under förmiddagen i dag har vi en fråga på föredragningslistan som kommer att få långtgående effekter för den gemensamma fiskeripolitikens framtid i Europa : att stärka dialogen med fiskeindustrin om den gemensamma europeiska fiskeripolitiken .
Inom Europaparlamentet har vi redan i flera år fört en dialog med fiskeindustrin .
Våra delegationer besöker också Europas fiskeregioner för att ställa frågor lokalt .
På så vis kan vi få en bättre inblick i problemen för dem som på ort och ställe dagligen måste leva och arbeta med de europeiska förordningarna .
Denna vecka besökte jag den s.k. gröna veckan , jordbruksmässan i Berlin , och jag hade där en diskussion med företrädarna för den tyska fiskerinäringen .
Frågan är högaktuell och explosiv , i synnerhet som vi står inför en reform av den europeiska gemensamma fiskeripolitiken år 2002 .
Principiellt skall politiken se till att alla intressen blir rimligt beaktade , och att det framför allt sker ett hållbart utnyttjande av fiskresurserna .
Kommunikationen mellan fiskerinäringen och gemenskapens organ måste löpa i båda riktningarna .
Industrin måste formulera sina behov och meddela kommissionen dem .
Å andra sidan måste kommissionen förbereda föreskrifterna och besluten och informera om dem .
Det som efterfrågas är en dialog , och inte en monolog .
Det har kommissionen insett .
Och endast om man har kännedom om problematiken , svårigheterna och möjligheterna till lösningar , vilka de berörda parterna bäst känner till , kommer man i framtiden att kunna fatta lämpliga beslut .
För att uppnå detta mål har kommissionen tagit två steg .
Med föreliggande förslag till förordning siktar kommissionen på att stärka de europeiska yrkesorganisationerna - med all rätt .
En dialog kan dock bara föras om ifrågavarande samtalspartner inom fiskerinäringen också får ekonomiskt stöd för att över huvud taget kunna delta i samtalen i Bryssel , dock utan att deras oberoende undergrävs .
För detta har ca 400 000 euro avsatts i år .
Huruvida dialogen blir framgångsrik kommer dock enbart att bero av hur kommissionen i de lokala regionerna kommer att kunna göra de komplexa tekniska aspekterna förståeliga med hjälp av sina informationsåtgärder .
Jag stöder därför uttryckligen dagens initiativ från kommissionen .
Samtidigt måste jag ändå uttala ett stort " men " .
Det gäller nämligen det andra steget , som Miguélez också har nämnt här .
Det handlar om reformen av den viktiga rådgivande kommittén för fiske och vattenbruk .
Detta är grunden för dialogen .
Varför rådfrågades inte Europaparlamentet när det gällde utformningen , organisationen och uppgifterna för detta så viktiga mellanled i den eftersträvade dialogen , dvs. just den rådgivande kommittén för fiske och vattenbruk ?
Detta är en brist , som vi kommer att fortsätta att kritisera .
Ytterligare några små " men " ser jag i svårigheterna att finna verkliga representativa företrädare för de olika sektorerna i den splittrade struktur som fisket utgör , med den geografiska mångsidigheten och den svaga organisationsstrukturen .
Här gäller det att äntligen skapa tillämpningsbara villkor .
Men förutsättningen är också att vi kanske överväger en ny organisationsstruktur inom fiskerinäringen .
Detta förutsätter dock återigen ett förtroende från de berörda yrkesfiskarna för politiken i allmänhet och för den europeiska gemensamma fiskeripolitiken i synnerhet .
Därför - det ber jag er - bör vi i framtiden göra så intensiva ansträngningar som möjligt .
Herr talman !
I går debatterade vi Cunhabetänkandet .
En av invändningarna från Europaparlamentets nederländska ledamöter var att de avtal som slutits i Nederländerna mellan staten och fiskerisektorn i syfte att på frivillig väg få avtal till stånd om efterlevnaden av fångstkvoten inte beaktas tillräckligt i detta förslag .
Om det är möjligt att få till stånd frivilliga avtal som har samma effekt som lagstiftning , i nära samråd mellan stat och samhällsorganisationer , då föredrar Arbetarpartiet sådana avtal framför onödig beskäftighet ovanifrån .
Det gäller naturligtvis även på Europanivå .
Jag är därför mycket nöjd med betänkandet av min kollega Miguélez Ramos .
Även om vi hade radikalt olika uppfattningar om Cunhabetänkandet stöder jag helhjärtat hennes förslag om att få en förstärkning av rådgivande kommittén för fiske till stånd .
Jag gratulerar henne till betänkandet .
Jag har i sammanhanget bara en randanmärkning .
Den rådgivande kommittén kan fungera väl endast om den är representativ för de olika sektorer som är involverade i fiskeripolitiken och om också unionens alla fiskerinationer är företrädda i kommittén .
Ännu så länge är det inte tal om detta .
Vår grupp kommer därför att rösta för ändringsförslag 3 , vilket syftar till att utöva ett visst tryck i den riktningen , och jag riktar också en uppmaning till Europeiska kommissionen att tillse att rådgivande kommittén är representativ , och att den även i fortsättningen kommer att vara beskaffad på det sätt som jag nyss beskrev .
Till sist , herr talman , kan jag meddela er att min grupp kommer att rösta för Miguélez Ramos resolution , eftersom denna ger ett viktigt bidrag till Europeiska unionens fiskeripolitik .
Herr talman !
Allt som kan stimulera och främja en dialog är värt att välkomna och en närmare dialog mellan fiske- och vattenbruksindustrin är något som måste uppmuntras .
Men inte bara industrin - vi måste utvidga dialogen till att omfatta organisationer som är aktiva på miljö- och utvecklingsområdet och låta specialiserade forskningsorgan få en mer framträdande roll .
Ett ömsesidigt kommunikationsflöde måste uppmuntras , inte bara envägskommunikation .
Mitt parti har alltid förespråkat ökat samråd med industrin .
En avgörande fördel med en regionalt förankrad strategi för den gemensamma fiskeripolitiken skulle vara att de direkt berörda , det vill säga fiskarna själva , tog del i beslut som påverkar dem .
Härigenom främjas målet att bevara fiskeresurserna genom ett hållbart fiske och de samhällen i Europa som är beroende av fisket erbjuds en långsiktig livskraft .
Utöver alla reformer från den rådgivande kommittén , vilka ingår i gemenskapens nuvarande utvärdering av den gemensamma fiskeripolitiken , har Europa en annan möjlighet att hitta bättre sätt att göra fiskarna delaktiga i genomförandet av fiskeriåtagandena , genom att utvidga regionaliseringsprincipen .
Genom att involvera industri och övriga berörda parter på orten skulle man skapa ett system som bättre avspeglar fiskeindustrins behov och främjar snarare än hindrar överensstämmelsen med den gemensamma fiskeripolitiken .
Genom att även säkerställa ett fungerande samråd med det civila samhället , i synnerhet fiskenäringen och miljöorganisationerna , säkerställer vi att gemenskapens fiskeripolitik korrekt avspeglar målen om bevarande av fiskeresurser och en hållbar utveckling inom fiskerisektorn .
Men de icke-statliga organisationernas deltagande måste vara meningsfullt , inte bara symboliskt , och vi måste arbeta hårt för att se till att så är fallet .
Att införliva dem som arbetar i fiskeindustrin i beslutsprocessen och stödja fiskarna är en nödvändig förutsättning för all framtida fiskeripolitik om den skall lyckas och en väsentlig del av den gemensamma fiskeripolitiken .
I går fanns meningsskiljaktigheter kring delar av Cunhabetänkandet , framför allt förslaget om sanktioner i form av minskade kvoter .
Skall samrådet vara meningsfullt är detta exakt den typ av förslag som vi måste rådfrågas om och jag beklagar att mitt förslag om att avsätta tid till detta inte gick igenom .
Jag hoppas att vi kan lära av misstagen och mena det när vi - som i detta betänkande som jag stöder - säger att vi vill förbättra kommunikationen och samarbetet med fiskeindustrin och de som berörs av fisket .
Herr talman !
Utan att höra de övriga EU-institutionerna har kommissionen inrättat en kommitté för fiske och vattenbruk .
Till samarbetspartner har kommissionen framför allt valt organisationer som är företrädda i gemenskapen .
Man vill inte att kommittén för fiske och vattenbruk är en talesman för nationella intressen .
Det är ändå precis vad den är .
Den är det åtminstone ur Finlands och Östersjöns synvinkel .
Medlemskapet i organisationen Europêche som är företrädd i gemenskapen är för dyrt för finländska fiskare .
De kan inte delta i organisationens verksamhet eftersom de inte har råd att betala medlemsavgifter .
Således försvaras inte deras intressen i de organisationer som kommissionen valt till sina samarbetspartner .
Fiskarna har inte råd med en representation i EU , men fiskodlarna har .
De är kapitalister inom fiskeribranschen .
Detta ställer gemenskapens fiskeripolitik i en egendomlig dager i vårt land .
Man lyssnar bara på fiskodlare , kapitalister , men inte på proletärer eller de fria yrkesutövare som på fria havsområden fångar fria fiskar , dvs. fiskarna .
Dessutom fiskar man hos oss i Norden även i insjöar , vilket man inte i EU tar hänsyn till .
Det här med de överstatliga organisationernas representativitet är en problematisk fråga eftersom EU inte i tillräcklig utsträckning fäster uppmärksamhet därvid .
Den överstatliga organisationen Europêche är ineffektiv .
Den är icke-representativ , dess beslut är inte bindande för medlemsorganisationerna , det är medlemsstaternas storlek och pengar som avgör , och som överstatliga intressen klassas där sådana frågor som i själva verket ligger i nationella intressen .
Komissionens viktiga uppgift är att tillämpa denna förordning , så att de organisationer som är företrädda i gemenskapen skall bli mera representativa , och att även sådana fiskare som inte har råd med medlemskap i en intresseorganisation på EU-nivå får sin röst hörd .
Herr talman !
Ledamöterna i Gruppen Union för nationernas Europa kan bara instämma med intentionerna i ett förslag till förordning som syftar till att stärka dialogen med de yrkesverksamma inom fiskerisektorn .
Men samtidigt måste vi säga att vissa av metoderna för att organisera dialogen är mycket förbryllande .
För det första behovet av att stärka dialogen .
Den gemensamma fiskeripolitiken omfattar Europeiska unionens samtliga aktörer , men den måste svara mot en mångfald av olika situationer , beroende på fiskezon , båtarnas hemmahamn , traditioner , de fiskeredskap som används , den lokala marknadsorganisationen , osv .
Detta till den grad att en del klarsynta människor har ställt sig frågan om en väl fungerande samordning av ländernas nationella politik inte skulle vara att föredra framför en enhetlig gemenskapspolitik .
Hur det nu än förhåller sig med det är dagens politik enhetlig och de yrkesverksammas situation mångskiftande .
Därför är det så mycket viktigare att organisera täta kontakter med de yrkesverksamma för att beakta deras behov och undanröja de perversa effekterna av vissa förordningar , eller undvika att man rätt och slätt avstår från att tillämpa dessa förordningar , vilket tyvärr ibland sker , eftersom de fullständigt saknar verklighetsförankring .
Detta är skälet till att ledamöterna i vår grupp kommer att rösta för de tre ändringsförslag som har lagts fram i dag .
Dessa syftar till att förbättra arbetet i den rådgivande kommittén för fiske och vattenbruk , knyta kommittén närmare till yrkesutövarna och medlemsstaternas behov , samt kräva att kommissionen lägger fram en årlig rapport för rådet och Europaparlamentet om överläggningarna i kommittén .
Samtliga gemenskapens institutioner , och inte bara kommissionen , är nämligen intresserade av denna diskussion , för att kunna bidra till att ge den gemensamma fiskeripolitiken en inriktning som överensstämmer med våra fiskeflottors legitima intresse .
Vissa inslag i reformen inger oss dock en djup känsla av olust , eftersom kommissionen låter påtryckningsgrupper av mycket skilda slag ta plats i den rådgivande kommittén .
Dessa är för övrigt till största delen hemmahörande i Bryssel och verksamma inom en mycket bred sfär - utveckling , miljö , konsumentfrågor osv .
På fiskarsidan vill kommissionen samtidigt , med hjälp av gemenskapsanslag , på bred front driva upp europeiska branschorganisationer som för närvarande bara existerar på papperet .
Det verkar som om kommissionen med hjälp av en mängd olika deltagare försöker uppväga de nationella organisationerna , som likväl är organiserade , förankrade och fullt representativa .
Det hela ser ut som om kommissionen försöker undvika diskussioner med samtalspartners som är svåra att styra och helt utan underlag skapa en fogligare samverkansstruktur som exakt återspeglar den behagliga bild av kommissionen och dess idéer som kommissionen förväntar sig .
Än mer oroande är att man till slut undrar hur många andra sektorer som redan har organiserats på detta sätt och om det inte i Bryssel har upprättats ett vidsträckt nätverk av organisationer utan verklig representativitet , till största delen finansierade genom gemenskapsbidrag och som deltar i till stor del konstlade samråd .
Det exempel vi i dag undersöker ger oss anledning att tro att risken är stor att denna hypotes är sann .
Under dessa omständigheter skall institutionerna i Bryssel inte förvåna sig över att de förlorar kontakten med folkopinionen .
Medlemsstaterna borde se allvarligt på detta , om de inte vill att de nationella demokratier som de företräder snart skall se sig utmanövreras av konturlösa påtryckningsgrupper .
När det gäller den sektor som för stunden sysselsätter oss , nämligen fiskerinäringen , tycks det oss absolut nödvändigt att tillse att de olika aktörerna i den rådgivande kommittén är väl representativa .
Alla medlemsstater som berörs av fisket bör vara företrädda , liksom yrkesgrupperna i dessa .
Det är dessa grupper vi skall utgå ifrån , och inte konstlade organisationer .
Herr talman !
Det är positivt att kommissionen tar initiativ för att förstärka dialogen med fiskeriorganisationerna .
Kommissionen måste känna till vad som sker på gräsrotsnivå .
Vi har inget behov av en kommission som utfärdar regler utifrån ett elfenbenstorn .
Samråd med sektorerna är nödvändigt för att man inte skall utfärda regler som inte är möjliga att genomföra i praktiken .
Det är likaledes nödvändigt med en dialog för att få en klar bild av olika intressen för att kunna fatta väl avvägda beslut .
Med det nu föreliggande utkastet till förordning avser kommissionen att förstärka de europeiska yrkesorganisationerna .
Det finns säkert en del att säga om detta .
Såväl fiskerisektorn som kommissionen har intresse av förekomsten av en europeisk paraplyorganisation .
För fiskerisektorn är det en viktig plattform för att få kommissionen att ytterligare uppmärksamma de gemensamma problemen .
Och kommissionen vet bättre vad den har att rätta sig efter om sektorn talar med en röst .
Men vi får ändå inte glömma bort att fiskerisektorn i allra högsta grad är en sektor med nationella motsättningar .
Om man talar med en vanlig fiskare kommer man att upptäcka att det som han ser det inte finns några europeiska fiskare .
Den europeiska flottan består av belgiska fiskare , danska fiskare , nederländska fiskare och så vidare , och de är i stor utsträckning konkurrenter till varandra .
Genomsnittsfiskaren har också mer förtroende för sin nationella intresseorganisation än för en europeisk där funktionärerna huvudsakligen utgörs av företrädare från andra medlemsstater .
Denna realitet får vi inte glömma bort .
Vi får inte heller betrakta en europeisk organisation som en ersättning för nationella organisationer , utan som ett komplement .
Europeiska kommissionen bör också fortsätta att föra samtal med de nationella organisationerna .
Detta för mig in på det ändringsförslag som min grupp har lagt fram om den rådgivande kommittén .
Det är sant att kommissionen inte har bett oss om ett yttrande med avseende på sammansättningen av den kommittén .
Men kommissionen kommer förhoppningsvis inte att ta illa upp om jag oombedd ändå kommer med en rekommendation .
Den 16 juli 1999 gick kommissionen och näringslivet med på en kompromiss om den nya rådgivande kommittén .
De kom då överens om att alla unionens medlemsstater , försåvitt de är fiskerinationer , måste vara företrädda i denna .
Intressemotsättningar gör det som sagt omöjligt för olika medlemmar av yrkesförbunden att ge sitt mandat till någon av annan nationalitet .
Den rådgivande kommittén sammanträdde nyligen i ny sammansättning .
Men tyvärr måste jag konstatera att det inte blivit mycket av med den balans man kommit överens om .
I kommittén är vissa nationaliteter kraftigt överrepresenterade , medan ett antal andra medlemsstater inte alls är företrädda .
Det var faktiskt skäl nog för den förre ordföranden för den rådgivande kommittén , under vars ledning kompromissen kom till stånd , att vägra att leda kommitténs första sammanträde .
Europeiska kommissionen kommer kanske att invända att representativitet innebär mer än en rättvis fördelning över medlemsstaterna .
Naturligtvis är det också så .
Det måste också handla om en rättvis fördelning över sektorerna .
Men vad jag skulle vilja veta av kommissionen är följande : " Varför har ni inte hörsammat kompromissen från den 16 juli där det tydligt står att det också måste vara tal om en rättvis fördelning vad nationalitet beträffar ? "
Jag vill därför framföra en angelägen rekommendation med adress till kommissionen .
Ompröva sammansättningen av den nya rådgivande kommittén .
Om ni vill ha en god dialog med de berörda sektorerna , om ni lägger vikt vid att skapa stöd för er politik , se då till att vi får ett representativt förhandlingsorgan .
Herr talman !
Precis som mina kollegor har gjort och precis som det framkommer i Miguélezbetänkandet vill jag också kommentera kommissionens godtyckliga arbetssätt .
Det är absurt att varken parlamentet eller rådet rådfrågades innan man påbörjade omorganiseringen av den rådgivande kommittén för fiske och att man nu dryftar förslaget till förordning för att förstärka dialogen mellan kommissionen och sektorn .
Man rådfrågar med andra ord inte om den normgivande grunden men däremot om de kompletterande aspekterna .
Inte om de regler som skall gälla för dialogen utan om hur den redan inrättade dialogen skall förstärkas .
Dessutom har den omorganisering som kommissionen har genomfört av ett så viktigt organ som den rådgivande kommittén , det enda organ som finns där sektorn involveras i de beslut som berör den , väckt både stark kritik och tvivel såväl i parlamentet som i rådet och i sektorn själv , där man anser att en stor del av fiskerisektorn inte är tillräckligt företrädd .
När nu detta väl är sagt och för att inte bli långrandig , tack och lov för de ekonomiska medlen i förslaget .
Det återstår bara att tacka Miguélez för betänkandet samt försvara de ändringsförslag där man åläggs att till oss översända en årlig rapport om innehållet i de debatter som hålls i de arbetsgrupper som bevakar förordningen i fråga .
Jag välkomnar också den begäran som framkom i Gallaghers yttrande , å utskottets för industrifrågor , utrikeshandel , forskning och energi vägnar där man dessutom begär detaljerad information om fördelningen av fonder till de medlemsländer och föreningar som kan gynnas av förslaget .
Herr talman !
Jag skall fatta mig kort .
Jag stöder detta betänkande och gratulerar föredraganden till hennes arbete .
Socialistgruppen välkomnar kommissionens reform av den rådgivande kommittén för fiske , för att skapa en mer fruktbar ömsesidig dialog mellan kommissionen och industrin .
Vi välkomnar att nya sektorer av industrin och ett bredare urval av yrkeskårer införlivas i kommittén , i synnerhet inom vattenbruk och saluföring .
Vi välkomnar att antalet ledamöter i plenarkommittén begränsas till förmån för större effektivitet .
Vi känner alla till farorna med att öka antalet ledamöter på bekostnad av effektiviteten .
Kommissionen verkar ha beaktat detta .
Vi välkomnar att forskningsorganisationerna ges en mer framträdande roll och att fyra arbetsgrupper inrättas .
Den första skall ansvara för tillgången till resurser och förvaltningen av fiskeriverksamheten , den andra för vattenbruk , fisk , skaldjur och musslor , den tredje för marknader och handelspolitik och den fjärde för ekonomi och strukturella sektorsanalyser .
Vi är positiva till prioriteringen av organisationer på gemenskapsnivå i ett försök att undvika att debatten domineras av nationella intressen , men vi erkänner att en del nationella uppgifter måste inhämtas på lämplig nivå .
Vi kommer att stödja detta betänkande , och lovar samtidigt att vara fortsatt vaksamma för att säkerställa att de så lovande strukturella förändringarna omsätts i praktiken , och att den nya rådgivande kommittén för fiske och vattenbruk fungerar som ett effektivt språkrör för alla sektorer och alla delar av industrin .
Herr talman !
Det är kanske ovanligt att jag yttrar mig om detta förslag när jag inte är ledamot av fiskeriutskottet .
Å andra sidan företräder jag - särskilt i västra Skottland - ett mycket stort antal fiskare och deras familjer och utsatta samhällen som för sin existens är beroende av att Europeiska gemenskapens fiskeindustri fortsätter att gå bra , och av att gemenskapen är uppmärksam på de utsatta och ofta avlägsna regioner i gemenskapen som är mest beroende av den .
Det är mycket lovvärt att säga att rådgivande kommittén för fiske inte bara skall vara en mötesplats för nationella intressen , särskilt om nationella intressen enbart tolkas som medlemsstaternas intressen , i enlighet med de proportionalitetsprinciper som styr medlemsstaternas representation i gemenskapens organ .
Det finns en annan princip som skulle vara proportionerlig i förhållande till det arbete som uträttas inom industrin och förvisso i förhållande till andelen fiskevatten och kuststräckor som olika regioner av gemenskapen bidrar med .
Jag ber ledamöterna göra ett litet experiment .
Tänk er att Skottland utesluts ur gemenskapen .
Hur mycket fiskeindustri skulle då bli kvar ?
Fundera nu över följande fråga .
Hur effektivt är den skotska fiskeindustrins röst företrädd i gemenskapens institutioner , så som de ser ut i dagsläget ?
Svaret är : alls inte särskilt effektivt !
Därför skulle det verkligen vara en god sak om detta betänkande kunde åstadkomma att fiskarna , miljöintressena och det civila samhällets övriga intressen företräddes långt mer effektivt .
Några stora framsteg tror jag inte vi gör genom detta betänkande , men något litet vore välkommet .
Herr talman , fru kommissionär , ärade kollegor !
Jag vill börja mitt anförande med att tacka föredragande Miguélez för ett väl genomfört arbete när det gäller en fråga av så stor vikt och social återverkan som en förstärkning av dialogen mellan kommissionen och den berörda sektorn har vid tillämpningen av den gemensamma fiskeripolitiken .
Föredraganden säger , vilket jag också menar , att det är ganska märkligt att kommissionen rådfrågar parlamentet i frågor som vi kan betrakta som sekundära för utformningen av dialogen och att man inte har hänskjutit frågan om sammansättning , organisation och verksamhet för den rådgivande kommittén för fiske , det egentliga forumet när det gäller att anordna dialogen , till parlamentet .
Jag menar att Europaparlamentet , som medborgarnas direkta och demokratiskt valda företrädare , borde ha uttalat sig om myndigheten i fråga och om representativiteten för de undersektorer som där ingår .
Nåväl , nu är det bara att vänta och se hur den nya kommittén kommer att fungera innan vi utvärderar verksamheten , vilket också är en anledning till att jag anser att det som sägs i Miguélez betänkandet beträffande den finansiella kontrollen av avgifterna och större öppenhet i förvaltningen , så att såväl parlamentet som rådet skall informeras så uttömmande som möjligt , så att vi alla gemensamt kan fullborda den förstärkning av dialogen som Europeiska kommissionen eftersträvar .
Jag hoppas att kommissionen noterar våra anmärkningar och vår oro , vi kommer nämligen att hålla oss väl informerade om utvecklingen av och verksamheten i den nya kommittén , med vilken vi från Europaparlamentets fiskeriutskott hoppas få ett gott samarbete , så att den sociala och sektoriella dialogen om fiske verkligen kan förstärkas .
Herr talman !
Som kristdemokrat skulle jag vilja göra en bedömning av kommissionens föreliggande förslag på två punkter .
Till att börja med respekteras subsidiaritetsprincipen , länderna är delaktiga på ett tillfredsställande sätt och för det andra beaktas organisationer eller lokala organisationer i tillräcklig utsträckning .
I den bemärkelsen är jag glad över att det skall bli en förstärkt rådgivande kommitté , som kanske också kan utöva mer inflytande på fiskeripolitiken .
Så långt är jag positiv .
I fråga om det verkliga innehållet är jag mindre positiv .
Jag konstaterar att förslaget på åtminstone två punkter är ett misslyckande .
Till att börja med är inte alla medlemsstater företrädda , och det anser jag vara mycket negativt , för vi erkänner i detta parlament även medlemsstaternas subsidiaritet .
Det innebär att medlemsstater med en viktig fiskerisektor inte får saknas .
Det andra är att när organisationer och lokala organisationer blir delaktiga i fiskeripolitiken måste detta ske på ett rättvist och bra sätt , varvid den geografiska spridningen är av stor vikt .
På den punkten är förslaget helt enkelt misslyckat .
Det är av den anledningen som jag tillsammans med andra kolleger , bland andra kollega van Dam , kräver att man ändå sörjer för att det skapas en rådgivande kommitté med en viktig roll , men att den är representativ för hela sektorn och för hela Europa .
Konkret innebär detta att alla unionens fiskerinationer bör vara företrädda i kommittén .
I den gamla rådgivande kommittén hade man uppnått samförstånd om detta mellan sektorn och kommissionen .
Att de aktuella förslagen som lagts fram av yrkesförbunden förbigår detta är som jag ser det , och även utifrån en kristdemokratisk syn , någonting negativt .
Herr talman !
Jag skulle vilja börja med att gratulera vår kollega Rosa Miguélez Ramos till hennes arbete .
Framför allt till den sansade analys betänkandet innehåller och för att hon har satt fingret på den ömma punkten eller rättare sagt , punkterna , för här finns två grundläggande frågor som redan har betonats av flera kolleger och som parlamentet måste notera .
Den första är vår förvåning , jag skulle vilja säga häpnad , över att parlamentet nu hörs om aspekter angående den rådgivande kommittén för fiske- och vattenbruk när det inte i tid hördes om dess sammansättning .
Förra året godkände kommissionen själv , som vi vet , beslut nr 478 / 99 som denna rådgivande kommitté hade skapat , och då hördes inte parlamentet i en så viktig fråga som den om fiskeorganisationernas representation och den viktiga roll som dessa har i utformningen och förvaltningen av den gemensamma politiken .
För mig är det obegripligt att parlamentet inte har hörts !
Det är ett rent mysterium .
Vissa förhållanden saknar skäl .
Jag vet inte om det finns några skäl till att parlamentet inte skulle höras som jag inte känner till .
Den andra anmärkningen är att vi hyser många betänkligheter angående representationen i dessa organ .
Exempelvis är inte ett land som mitt , Portugal , som är en fiskerination på europeisk nivå och som har den femte största fiskeflottan i unionen , företrätt på ett rättvisande sätt .
Jag är häpen , för mig är detta verkligen ett mysterium .
För att avsluta den andra frågan , det vill säga den andra ömma punkten , och med hänsyn till den rådgivande kommitténs luckor och representationen där , är det viktigt att avsätta och överväga finansiellt stöd till andra organisationer som inte ingår i den rådgivande kommittén .
Herr talman !
Jag välkomnar detta betänkande och tackar fru Ramos för hennes inledning som var lättfattlig och konstruktiv .
Det är meningsfullt med denna insats för att främja en bättre dialog mellan Europeiska unionen och de aktiva inom fisket .
I den del av Europeiska unionen som jag kommer från , en avlägsen region , har vi alltid haft särskilda svårigheter att vinna gehör för tanken om en gemensam fiskeripolitik hos fiskarna .
Eftersom MacCormick tog upp frågan - och jag har varit inne på den tidigare - är Irlands ställning besvärlig , för om Irland uteslöts ur Europeiska unionen skulle mycket fisk försvinna samtidigt .
Av tradition brukade irländska fiskare inte fånga den här fisken , eftersom det som en del av er vet under en period av vår historia i lag var förbjudet att ta upp fisk på irländska fartyg .
Detta förhållande levde till stor del kvar fram till början av 1900-talet och därför fiskade folk så sent som 20 år före vårt inträde i Europeiska unionen i gammalmodiga fiskebåtar .
Hur som helst är det ett faktum att fisk till ett värde av runt 700 miljoner euro - och kanske rentav mer , eftersom priset på fisk har ändrats - kommer från irländska fiskevatten .
Som ett resultat av att strukturfondsstödet till Irland har minskat i den ekonomiska tillväxtens spår , kommer värdet på den fisk som skulle fångas i irländska vatten om inte Europeiska unionen fanns om ett par år att överstiga det totala strukturfondsstöd som utbetalas till Irland .
Detta gör det ändå svårare att vinna gehör för förslaget .
Jag känner inte till att detta gäller något annat land i Europeiska unionen .
Skottland är en del av Förenade kungariket och får sin beskärda del tillsammans med Förenade kungariket , men Irland är det enda undantaget .
Det här mig veterligt den enda naturresurs som alla medlemsstater går med på att betrakta som Europeiska unionens gemensamma egendom .
Detta innebär inte att vi inte behöver fullfölja denna dialog .
Utvidgningen av tjugomilsgränsen , som parlamentet har godkänt , kan vara en del av lösningen och bidra till att tillfredsställa lokala fiskare och ge dem större kontroll över sina liv .
Jag vill inte se någon ny nationalisering , men en regionalisering skulle förvisso vara till hjälp för Skottlands och Irlands problem .
Herr talman !
Jag skulle vilja inleda med att säga att de ofta förekommande ändringarna i lagstiftningen som rör den gemensamma fiskeripolitiken visar på den dynamik som finns på detta område .
En dynamik som inte kunde komma till uttryck inom ramen för funktionen av den föregående rådgivande kommittén för fiske , och det var därför detta lagstiftningsförslag lades fram .
Målet med detta förslag är att skapa en effektivare och mer påtaglig relation mellan kommissionen och den rådgivande kommittén för fiske .
Det krävdes tre års arbete för att kommissionen skulle komma fram till detta förslag .
1997 fick en oberoende byrå i uppdrag att genomföra en undersökning , och den ledde till två slutsatser .
Den första är att fiskeripolitiken inte är av intresse enbart för fiskeindustrin utan att den nu även berör andra delar av samhället .
Och det är någonting som vi måste beakta .
För det andra svarade inte det sätt som den rådgivande kommittén fungerade på mot de behov som hanteringen av komplicerade frågor krävde .
Nå , lagstiftningsförslaget består av tre delar : Den första gäller reformen av den rådgivande kommittén , som nu består av 20 medlemmar , i stället för 45 , och vars deltagare till 60 procent kommer från fiskeorganisationerna , till 25 procent från industri- och affärsföretagen i branschen och till 15 procent från miljöorganisationerna .
Man har alltså försökt ordna det så att kommissionen skall kunna inhämta åsikter inte bara från yrkes- och branschfolket utan även från själva samhället .
Lagstiftningsförslagets andra del gäller åtgärder för att stärka de organisationer som företräder de kretsar som berörs av den gemensamma fiskeripolitiken , särskilt de europeiska yrkesfiskarorganisationerna .
Den tredje delen handlar om att förbättra kontakterna mellan Generaldirektoratet för fiske och dessa kretsar .
Lagstiftningsförslaget handlar om de två sistnämnda punkterna , men jag vill upprepa att det slutgiltiga förslaget föregicks av en lång period av överläggningar avseende kommitténs sammansättning .
Den 26 oktober var detta förslag föremål för en första granskning i rådet , som redan väntar på parlamentets yttrande för att kunna gå vidare i sitt arbete .
Jag vill särskilt ge komplimanger till Ramos för den enastående kvaliteten på hennes betänkande , liksom jag vill ge komplimanger till parlamentets fiskeriutskott för vårt mycket goda samarbete och för arbetet med denna text .
Jag skulle vilja kommentera ändringsförslagen och redogöra för kommissionens ståndpunkter .
Parlamentets utskott har utarbetat tre ändringsförslag .
I det första tar man upp parlamentets önskan om att yrkesorganisationernas betalningar skall kontrolleras noga , så att de exakt motsvarar de mål som har fastställts i lagstiftningsförslaget .
Kommissionen instämmer i detta och godkänner ändringsförslaget .
Vad beträffar det andra ändringsförslaget , instämmer kommissionen i parlamentets åsikt att all information om kommitténs arbete och om de många kontakter som kommittén har måste redovisas .
Att sammanställa en årsrapport är , med tanke på verksamhetens omfång , ett mycket krävande arbete för det redan tungt belastade generaldirektoratet för fiske , som inte skulle medföra några tydligt urskillningsbara vinster .
I det tredje ändringsförslaget inbegrips innehållet i det andra , och det handlar om representationen i den rådgivande kommittén , det vill säga om deltagande av alla nationaliteter .
Vi håller med om att det bör säkerställas att hela sektorn på ett balanserat sätt företräds i kommittén , men vi tvivlar på i vilken utsträckning - och det har framkommit såväl i undersökningarna som under dialogen - denna balans bör fastställas på grundval av nationalitet .
Kommissionen vill stärka de europeiska organisationerna , som har alla möjligheter att själva ombesörja den nationella representationen eller representationen för särskilda kategorier , när de bedömer att det är nödvändigt .
Jag skall avsluta med att säga att kommissionen godtar ändringsförslag 1 , i vilket gemenskapen uppmanas att stärka den offentliga kontrollen , men att den anser det vara lämpligt , av de skäl som jag har redogjort för ovan , att förkasta ändringsförslagen 2 och 3 .
Tack så mycket , fru kommissionär .
Herr talman !
Jag skulle vilja ställa en fråga till kommissionären .
Jag tror att alla de ledamöter som har talat har ställt samma fråga till kommissionen .
Varför rådfrågade kommissionen inte parlamentet om reformen av den rådgivande kommittén när parlamentet under den föregående mandatperioden , när förslaget fortfarande låg på bordet , begärde detta ?
Jag skulle vilja att kommissionären besvarade den här frågan men framför allt att hon formellt går i god för att detta inte kommer att upprepas . .
( EL ) Herr talman !
Frågan är förståelig , men jag vill upprepa att kommissionen arbetar med fördraget som grund och inom en bestämd ram , som den måste respektera .
Denna kommitté är en gemenskapskommitté , och ingenstans finns det föreskrifter om samråd med parlamentet vid reformeringar av denna slags kommittéer , vilka upprättas av kommissionen .
Herr talman !
Innan vi övergår till omröstning skulle jag gärna vilja få en liten verifiering .
Så sent som en kort stund före det att vi inledde detta sammanträde fanns det fortfarande ingen definitiv röstningslista tillgänglig .
Jag skulle gärna vilja att ni bekräftade det som vi redan fått höra av funktionärerna , nämligen att omröstning med namnupprop gäller för ändringsförslag 3 .
Jag vill i samband med ändringsförslag 3 också anmärka att det inte bara är författat av EDD-gruppen , utan även av ett tiotal andra ledamöter från PPE-DE-gruppen .
Ja , ledamot van Dam .
Omröstningen med namnupprop har tagits med i beräkningen .
Jag förklarar debatten avslutad .
Omröstning kommer att äga rum .
( Parlamentet antog lagstiftningsresolutionen . )
Röstförklaringar Herr talman !
Är det inte en aning sadistiskt av oss att alltid diskutera fiskerifrågor på fredagar , när fisken hos oss hamnar i stekpannan ?
I Camogli , nära Genua , min födelsestad , finns det en enorm stekpanna där man varje år steker fisk som sedan delas ut gratis till stadens invånare .
Detta säger jag för att förklarar varför jag är intresserad av fiskerifrågor och varför jag röstade för den här resolutionen .
Det är rätt att medborgarna tillfrågas och , även om kommissionär Diamantopoulou just har förklarat för oss att kommissionen inte behöver fråga medborgarna , så skulle jag vilja föreslå att man vid utfrågningar i ämnet även ger tillträde åt de äldre fiskarna . - ( PT ) Jag röstade emot såväl i slutomröstningen som angående lagstiftningsresolutionen , eftersom en majoritet i parlamentet tyvärr inte , kanske för att den lydigt lyssnade på den muntliga opposition den närvarande kommissionären uttryckte i debatten , godkände ändringsförslag 3 som Gruppen för demokratiernas och mångfaldens Europa och andra ledamöter individuellt hade ingivit .
Det går inte att förstå resultatet , eftersom kritiken mot kommissionen i samma debatt för att den inte rådgjorde med parlamentet om reformen av sammansättningen av den rådgivande kommittén för fiske var praktiskt taget generell .
Just ändringsförslag 3 var det enda som grep in på det här planet på ett oumbärligt sätt för att garantera en verklig representation i denna partnerstruktur , och övervinna dess obalanserade och mycket fiktiva karaktär .
Det är beklagligt att till och med i en så här enkel fråga fortsätter den gemensamma fiskeripolitiken att fungera på ett dåligt sätt .
 
Biståndsarbetare i Colombia Nästa punkt på föredragningslistan är debatten om följande muntliga frågor till kommissionen : B5-0006 / 2000 av Sauquillo Pérez del Arco för PSE-gruppen om skydd för biståndsarbetare .
B5-0007 / 2000 av Kreissl-Dörfler , Lipietz och Nogueira Román för ARE / EDN-gruppen om skydd för biståndsarbetare i Colombia .
Herr talman !
Jag vill inte vara dramatisk och jag vet att många ur civilbefolkningen utsätts för våld vid väpnade konflikter i olika länder .
Mellan 1992 och 1997 mördades emellertid 131 hjälparbetare , humanitär personal i FN : s tjänst som kämpar för de mänskliga rättigheterna på platser där konflikt råder .
Mellan den 1 januari 1994 och den 17 mars 1997 kidnappades vid 35 tillfällen 119 personer , alla hjälparbetare och humanitär personal .
1992 dog en FN-representant varje månad en våldsam död .
1993 dog en varannan vecka och 1994 en varje vecka .
Under de första två månaderna 1997 dog 9 samarbetspartner .
1996 utsattes 153 ombud från Röda korsets internationella kommitté för olika incidenter , inklusive mord och kidnappning .
Jag vill särskild påminna om de tre mördade läkarna från organisationen Läkare utan gränser - Spanien i Rwanda 1997 .
Nåväl , som vi säger i kompromissresolutionen , med vilken vi vill avsluta den här debatten , så är morden på samarbetspartnerna Iñigo Eguiluz och Jorge Luis Mazo från organisationen Fred och tredje världen den 18 november i Quibdó , 500 km norr om Bogotá vid Atratofloden , bara det sista i en lång rad av attentat .
Attentat inte bara mot personernas integritet utan mot de mänskliga rättigheterna , de internationella mänskliga rättigheterna och rätten för konflikternas offer att få hjälp , att förövarna döms samt att erforderliga åtgärder vidtas för att förhindra att den här typen av brott förblir straffria .
Den osäkerhet som biståndsarbetarna känner beror givetvis på att antalet väpnade konflikter har ökat , men även på att hjälporganisationerna är fler och att konflikterna i sig är av annan karaktär .
Det är inte längre fråga om konflikter mellan den reguljära krigsmakten , som kontrolleras politiskt , och några hierarkiskt styrda paramilitära rörelser med en tydligt angiven ideologi , där parterna i konflikten på ett eller annat sätt var ansvariga för hjälparbetarnas skydd , vars aktiviteter gynnade befolkningen .
I dag finns inte detta längre .
Hjälparbetarna och aktivisterna utsätts för stråtröveri .
Civilbefolkningen betraktas bara som en faktor till i konflikten , en del av såväl den politiska som militära strategin .
De humanitära aktiviteterna hindrar därför parterna i konflikten att nå sina mål , vilka ofta av etniska , religiösa eller kulturella skäl består i att eliminera en del av civilbefolkningen .
Inför en sådan verklighet är biståndsarbetarnas säkerhet en fråga med stor räckvidd som oroar parlamentet och som borde oroa såväl kommissionen , som finansierar mer än 180 icke-statliga organisationer i konfliktområdena , som rådet , som förtvivlat försöker bedriva en utrikespolitik i överensstämmelse med fördragen med främjandet av de mänskliga rättigheterna och med den säkerhetspolitik som just nu konkretiseras i humanitära gärningar .
Vi i parlamentet vill därför uppmana övriga institutioner att också känna oro .
Kommissionen genom att utforma ett meddelande om säkerhetsvillkoren för hjälp- och biståndsarbetare och genom att vidta åtgärder som kan garantera våra biståndsarbetares säkerhet .
Innan vi kommer till de åtgärder som föreslås av en del regeringar , som till exempel ett militärt skydd för biståndsarbetarna , måste vi lägga fram andra effektivare förslag .
Rådet kan genom GUSP främja de internationella mänskliga rättigheterna och en europeisk civil fredsstyrka kan kanske inrättas .
1999 firade vi femtioårsdagen av Genèvekonventionen för de mänskliga rättigheterna , den konvention som skyddar civilbefolkningen i väpnade konflikter och garanterar ett internationellt bistånd .
Det är ett instrument som är juridiskt förpliktande för alla länder och ändå blir det systematiskt förbigått .
Vi uppmanar rådets generalsekreterare att använda sig av Europeiska unionens begynnande kapacitet och främja de här principerna utanför Europeiska unionen .
FN : s generalsekreterare uppmanade i dagarna Säkerhetsrådet att genomdriva de internationella mänskliga rättigheterna genom att tillämpa kapitel 5 , 6 och 7 i Förenta nationernas stadga .
I dag ber vi er bara att bli mera medvetna och vidta åtgärder så att vi kan ta itu med ett problem som inte bara berör icke-statliga organisationer utan också grunden till vår uppfattning om världsordningen . .
( EL ) Kommissionen beklagar särskilt den tragiska händelsen , som är en av de som äger rum dagligen runt om i världen och som ledamoten också gav exempel på .
Kommissionen uttrycker sitt beklagande och betonar samtidigt ännu en gång det mod och det engagemang som visas av den humanitära personal som arbetar i dessa så farliga områden runt om i världen .
Särskilt när det gäller Colombia har kommissionens vid upprepade tillfällen för myndigheterna i Colombia betonat sin oro över denna fråga .
Vi fortsätter att övervaka situationen , och vi samarbetar kontinuerligt med medlemsstaternas ambassader i Bogotá .
Vad beträffar morden på Iñigo Eguiluz , som arbetade med ECHO-projekt , och prästen , har kommissionen och medlemsstaterna tryckt på de colombianska myndigheterna att genomföra undersökningar om detta brott .
Europeiska kommissionen och Spaniens ambassadör har träffat den colombianske vicepresidenten och insisterat på att de skyldiga till brottet måste ställas inför rätta .
Att rädda och skydda liv under dessa extraordinära omständigheter utgör en oskiljaktig del av den humanitära rätten .
ECHO : s roll i Colombia , och i andra länder , är att övervaka den humanitära situationen i landet , men även , särskilt i Colombia , att övervaka situationen för de människor som tvångsförflyttas , och det görs oavbrutna ansträngningar för att kontrollera att den humanitära rätten tillämpas .
Ledamoten underströk emellertid behovet av särskilda åtgärder från kommissionens sida för att garantera säkerheten för denna personal .
Ni hänvisade till ett redan existerande kommissionsdokument som är ett dokument om biståndspersonalens säkerhet från i maj 1998 i vilket prioriteringarna redovisas och de konkreta åtgärderna tas upp .
På grund av den förvärrade situationen , anordnade i april 1999 kommissionens kontor för humanitärt bistånd , ECHO ett seminarium om säkerhetsfrågor i Bogotá med Röda korsets internationella kommitté , och alla organisationer som är verksamma i Colombia uppmanades då att utarbeta en säkerhetsstadga och att i förväg meddela sina resor till Röda korsets internationella kommitté .
Detta för att säkerställa att de olika väpnade grupperna blir informerade om uppdragens humanitära karaktär .
Jag måste även betona att det förutom behovet av planering , åtgärder och personalutbildning även finns ett behov av finansiering .
Det är inte gratis att genomföra den humanitära hjälpen .
Av den anledningen inte bara uppmuntrar kommissionen det praktiska genomförandet av den humanitära hjälpen , utan den finansierar också verksamhet som avser att ge de personer som deltar i dessa uppdra en ökad kunskap och ett ökat medvetande om farorna .
Tillåt mig att ta upp några exempel på nya och tidigare initiativ som har tagits i detta syfte : Utarbetandet av dokumenten om den humanitära hjälpen , seminariet om säkerhet med partner i Lissabon , arbetsgruppen för personal i Bryssel om säkerhetsfrågor , införlivandet av frågorna om personalsäkerhet i ECHO : s handböcker samt sammanträdet för ECHO : s medarbetare , som kommer att äga rum i februari-mars i år av denna anledning .
Naturligtvis kommer Europaparlamentets förslag att beaktas , och eftersom det rör sig om en fråga som inbegriper mycket stora svårigheter och väldigt olika aspekter , är ett nära samarbete , de nya idéerna och förslagen mycket betydelsefulla även för kommissionens agerande .
Herr talman !
Mordet på biståndsarbetaren och missionären Iñigo Eguiluz och den colombianska prästen Jorge Luis Mazo vid Atratofloden i Colombia är en tragisk händelse och ännu en i raden av våldsamma dödsfall som de senaste åren har berört de volontärer som ägnar sina liv åt att uppnå fred och som dessutom förser de mest missgynnade med en kultur .
Det är därför logiskt att min grupp och parlamentet visar sitt deltagande och skickar ett kondoleansbrev till offrens familjer och ett budskap om stöd och hopp för de medarbetare som fortsätter med sitt arbete .
Samtidigt vill vi uppmana ansvariga institutioner att se till att lagen följs , och att kommissionen , rådets generalsekreterare och den colombianska regeringen gör vad som står i deras makt så att lag skipas och händelserna straffbeläggs enligt gällande lag .
Fängslandet av en förmodad brottsling är ett positivt tecken som vi lovordar , liksom vi lovordar president Pastranas vilja såsom den kom till uttryck vid hans senaste besök här i parlamentet .
Vi förstår svårigheterna , men vi vill ändå påminna regeringen om att stödet för Röda korset och FN : s flyktingorgan är något som alltid kan räkna med vårt stöd , liksom ansträngningarna av en rigorös tillämpning av 1998 års lagstiftning och föregående så att de här grupperna får ett rättsligt och reellt skydd .
Vi medger också att det är nödvändigt att förstärka de system som finns för att finna och rättsligt skydda biståndsarbetare och volontärer .
De arbetar i områden där konflikt råder , våldsamma och fattiga områden , områden där mörker råder och dit rättvisan inte når , därför måste vi försöka finna andra lösningar , andra typer av system .
Vi som lever i välfärd , de europeiska institutionerna och regeringarna , är bundna av en hederskodex och måste kringgärda dem som kämpar för de mänskliga rättigheterna med ett skyddsnät och fullständigt stödja rättvisan .
Medan vi försöker hjälpa till utifrån åstadkommer de fred och solidaritet inifrån , de tränger in i dunkla områden och ger hälsa och lösningar .
Det är den ädlaste versionen av ett tillmötesgående samhälle , vårt svar måste därför vara effektivt och ansvarsfullt .
Herr talman !
Kommissionär Diamantopoulous uttalande lugnar oss såtillvida att kommissionen är medveten om de problem som uppstår tack vare den bristande säkerheten för biståndsarbetare i vissa länder .
Sauquillo betonade såväl i sin muntliga fråga som i den redogörelse hon just lämnat att problemet inte är specifikt för ett visst land .
Det är sant att Colombia är ett av de länder som inte kan garantera biståndsarbetarnas säkerhet .
Det är dock inte bara Colombia det är frågan om .
Samma problem finns i många länder i Afrika och Asien , samt i andra områden .
I resolutionsförslaget uppmanas kommissionen att uttala sig i frågan .
Jag vet inte om det är det lämpligaste instrumentet , men det verkar som om kommissionen är beredd att arbeta i den här riktningen , och då är det förmodligen fördelaktigt om man började tänka på att utforma något slags dokument .
Det som enligt min mening inte verkar vara så meningsfullt är att öronmärka Colombia eller att stödja några av de ändringsförslag som lagts fram och där man till exempel föreslår att samarbetet skall brytas .
Stoppas samarbetet med sådana här länder kommer medborgarna att åsamkas stor skada .
Låt oss inte hindra detta samarbete , det är nämligen ett osjälviskt samarbete av människor som vet vilka risker de utsätter sig för .
Säger man å andra sidan att man kan vara utan ett regeringssamarbete så känner man inte till verkligheten .
Jag har besökt ett flertal områden i Colombia och förutom de normala faktorerna - det är ett svårt land - så finns ytterligare ett problem eftersom det finns olika grupperingar och man vet inte vilken av dem som kan mörda .
Utan regeringshjälp blir samarbetet absolut omöjligt .
Jag menar att debatten är viktig när det gäller att påminna kommissionen om vad som håller på att hända .
Kommissionen har lugnat oss med att säga att det är en fråga som oroar , men vi måste se situationen som den är .
Det internationella samarbetet måste fortsätta .
Europeiska gemenskapen måste fortsätta att föregå med gott exempel och visa vad ett internationellt samarbete är , vi måste stödja våra biståndsarbetare och det vore önskvärt att man härifrån , från gemenskapsinstitutionerna , medlemsländernas regeringar och givetvis mottagarländernas regeringar , garanterar säkerheten för de här människorna .
Först med ett förebyggande skydd .
Sedan med rättsliga åtgärder .
De colombianska myndigheterna försäkrar mig att ett rättsligt förfarande har inletts och att en person har häktats .
I Colombia är den dömande makten mycket självständig och den verkställande makten har ingen befogenhet att sätta sig över brottslighet utan man måste följa vanliga straffrättsliga förfaranden .
Kommissionär Diamantopoulou , jag uppmanar er att fortsätta på den väg ni har slagit in och jag hoppas att vi kan förbättra säkerheten för våra biståndsarbetare .
Herr talman !
Jag talar i dag som företrädare för de kolleger som står bakom det andra förslaget på dagordningen , som har förelagts parlamentet .
De beklagar att de inte kan närvara själva .
Även om jag inte är lika insatt i frågan är jag glad över detta tillfälle att företräda dem och Gruppen De gröna / Europeiska fria alliansen .
Som parlamentariker gör vi oss ofta skyldiga till klagomål på olägenheter i vårt liv , när vi reser mellan två , tre eller fyra städer , sitter på trånga kontor och så vidare .
Därför är det ett ögonblick som manar till ödmjukhet att inför parlamentet tala om detta ämne och begrunda de problem och faror som möter de modiga människor som ger sig ut som biståndsarbetare i tredje världen .
Vi kan bara stanna upp och tänka på förhållanden under vilka de lever , och tyvärr ibland också dör .
Med det vill jag ha sagt att min grupp och jag är besvikna över att våra kolleger i socialistpartiet enligt vårt förmenande tycks tappa bort behovet att fokusera på Colombia - även om de har rätt i att detta är ett generellt problem .
Det är viktigt att komma ihåg att president Pastrana besökte parlamentet så sent som i oktober och utfäste garantier om värnandet om de mänskliga rättigheterna , brottsbekämpning och upplösning av de paramilitära grupperna .
Dessa garantier har visat sig vara närmast värdelösa .
Vad som har gjorts är otillräckligt .
Enligt förslaget från min grupp måste kommissionen villkora sin närvaro och sitt arbete i landet genom att kräva en skärpning av lagarna rörande skydd av fördrivna arbetare och kräva att den colombianska regeringen garanterar deras fysiska säkerhet och materiella välbefinnande .
Det är riktigt att kommissionen måste vidhålla dessa krav .
I nästa stycke i förslaget står det att vi motsätter oss fortsatt stöd till den colombianska regeringen .
Men inte till det colombianska folket , eftersom det i nästa stycke står att vi bör fortsätta att ge stöd genom andra kanaler och styra stödet så att vi försäkrar oss om att de paramilitära grupperna inte får del av det , och att lag och ordning så snart som möjligt återupprättas i Colombia .
Hjälparbetarna är en besvärlig del av problemet , men inte hela problemet .
Det enda sättet att hejda dödandet är att upplösa de paramilitära grupperna och förse hjälparbetarna med lämpliga livvakter .
ECHO och kommissionen måste sätta press på regeringarna för att åstadkomma detta .
Herr talman !
Den 26 oktober förra året talade Colombias president , Pastrana , här i Europaparlamentet .
Han sade sig då vilja arbeta för mänskliga rättigheter i sitt land , för att de aktivister som arbetar med frågor som rör mänskliga rättigheter skulle få skydd , och för att skyldiga till mord och våldsbrott som främst begås av paramilitära grupper inte skulle få straffrihet , utan ställas till ansvar .
Mindre än en månad senare skedde de mord som är bakgrunden till dagens debatt .
En paramilitärgrupp angrep organisationen Fred och tredje världen , en organisation som med stöd av ECHO-programmet arbetar för humanitärt stöd till fördrivna jordbrukare .
En colombiansk präst och en spansk hjälparbetare dödades .
Den spanska hjälparbetaren arbetade för de fredsbrigader som med sin närvaro skall skydda aktivister för mänskliga rättigheter mot våld .
Dessa mord är bara några i den långa raden av övergrepp i Colombia , men denna gång dödades också en medborgare från ett EU-land .
Mord och försvinnanden tillhör den colombianska vardagen .
Exempelvis försvann helt nyligen två framstående talespersoner för bonderörelsen , bortförda av en paramilitär grupp , och de är inte återfunna .
Bakom större delen av denna terror står paramilitära grupper med mer eller mindre uppenbar koppling till landets egen militär och maktstruktur .
Upprepade gånger har det bevisats hur landets militär har varit direkt inblandad i olika våldsdåd .
Offren är civilbefolkning i områden där gerillan har stöd , den politiska vänstern , fackliga aktivister och de som arbetar för mänskliga rättigheter .
Den lagliga vänstern i landet har drabbats hårt .
Tusentals av dess företrädare , inklusive borgmästare och parlamentariker , har helt enkelt mördats .
Mycket sällan har förövarna straffats .
I ett sådant land är det inte märkligt att många söker sig till gerillan och till den väpnade kampen .
Det skall dock understrykas att även gerillan gör sig skyldig till våldsdåd som omöjligen kan försvaras .
Att uppnå en bättre respekt för mänskliga rättigheter i Colombia är helt avgörande för att det skall kunna bli en fredlig lösning på inbördeskriget i landet .
Fredsansträngningarna måste stödjas , samtidigt som den colombianska regeringen måste stå under ständig press , inte minst från Europeiska unionen vad avser mänskliga rättigheter .
Utländsk , dvs. amerikansk , militär inblandning måste avvisas .
Vår grupp , GUE / NGL-gruppen , har inte kunnat skriva under den kompromissresolution som har förhandlats fram .
Vi menar att den är helt otillräcklig i kritiken mot den colombianska regeringen .
Det är märkligt att man i punkt D i resolutionen berör en ockupation av ett Röda kors-kontor av jordbrukare , samtidigt som man inte på ett tydligt sätt tar upp de tusentals politiska mord som har skett i Colombia .
Vi har lagt fram två ändringsförslag tillsammans med Gruppen De gröna .
I det första ändringsförslaget vill vi att hjälp till den colombianska regeringen skall göras beroende av respekt för mänskliga rättigheter och att man skyddar dem som arbetar med dessa frågor .
I det andra ändringsförslaget vill vi utöka den humanitära hjälpen genom organisationer som är oberoende från Colombias regering , t.ex. de civila fredskårerna .
Om dessa ändringsförslag antas , blir denna resolution något bättre och tydligare .
Herr talman !
Bildandet av Röda Korset efter slaget vid Solferino var ett svar på en dittills okänd dimension av grymhet , det s.k. moderna totala kriget , som på ett avgörande sätt präglade 1900-talet .
Men i början av 2000-talet upplever vi en allt starkare utbredning av nya slags krig , i form av etniska konflikter i milis som stöter ihop , parter i ett inbördeskrig , eller helt enkelt kriminella gäng .
Regeringarna är antingen inblandade , eller också är de helt eller delvis maktlösa .
Detta äventyrar naturligtvis också i stor utsträckning den humanitära hjälpen och utvecklingsstödet .
Därför är det vår uppgift inom Europaparlamentet att intensivt ägna oss åt denna fråga , att uppskatta vad människor inom utvecklingsstödet och inom den humanitära hjälpen här gör , men också se till att deras levnads- och arbetsvillkor förbättras .
Jag tror att vi här har mycket att ta igen .
Vi måste se till att Europeiska unionen också faktiskt lämnar hjälp överallt där exempelvis de icke-statliga organisationerna gör det på ett förebildligt sätt .
Vi har inte bara den problematiken i Sydamerika , utan denna vecka hade vi en debatt om Tjetjenien , för någon tid sedan en om Centralasien , och sedan hörde vi kollegan Madelin om Afghanistan .
Och alltid samma fenomen : Man drar tillbaka den humanitära hjälpen , eftersom ingen säkerhet kan garanteras .
Vissa icke-statliga organisationer visar på hur man ändå , med stora risker , kan lämna hjälp .
Men Europeiska unionen och även andra stora organisationer , exempelvis Röda korset , befinner sig alltför ofta på återtåg .
Vi måste se upp så att denna tendens inte fortsätter , ty den utnyttjas skamlöst av vissa regeringar , som säger att man vill lämna hjälp till respektive regering och inte direkt via de icke-statliga organisationerna på platsen .
Det är farligt , ty dessa regeringar utgör ju inte lösningar på problemet , utan är en del av problemet , och de är också orsaken till det .
Därför måste vi här verkligen se till att vi håller i trådarna även i fortsättningen .
Av den anledningen börjar vi som parlament att bli mycket besvikna på vår ansvarige kommissionär Nielsen .
Fru kommissionär , jag ber er också meddela kommissionären detta .
Missnöjet har under flera veckor tilltagit här i kammaren .
Vi hade administrativ kritik beträffande Bonino .
Men Bonino var närvarande .
Hon var inte bara närvarande i parlamentet , utan också i krisområdena .
Europeiska unionen hade ett ansikte när det gällde den humanitära hjälpen och utvecklingsstödet .
Här har kommissionen mycket att ta igen .
Vi börjar här långsamt - det hör jag i alla grupper - att utveckla en mycket kritisk hållning .
Jag anser att man i tid bör övergå till att återigen skapa gemensamma initiativ för att stabilisera den politiska miljön , stödja de icke-statliga organisationerna men också se till att Europeiska unionen är närvarande på platsen , där så krävs . .
( EL ) Herr talman !
Dialogen om så svåra frågor som den humanitära hjälpen , förvaltningen av den humanitära hjälpen och personalens säkerhet runt om i världen är verkligen mycket viktig , och Europaparlamentets roll är mycket betydelsefull .
Jag skulle dock vilja , det var därför som jag begärde ordet , säga några ord om kommentarerna om kommissionär Nielsen .
För det första närvarar han inte i dag på grund av att han befinner sig på resa i Sydafrika , för det andra har han under dessa tre månader verkligen besökt många krishärdar och för det tredje har arbetat hårt , och han har redan lagt fram förslag till kommissionen både om en fullständig omstrukturering av och om nya förordningar om förvaltningen av den humanitära hjälpen och om nya former av samarbete med de icke-statliga organisationerna .
Jag förstår och instämmer med många av ledamöternas kommentarer om de problem som finns , men jag tycker att det är överdrivet att en kommissionär som har varit kommissionär i tre månader och som redan har uträttat viktigt arbete kritiseras så hårt .
Tack så mycket , Diamantopoulou .
Jag har mottagit fyra resolutionsförslag i enlighet med punkt 5 , artikel 42 i arbetsordningen för att avsluta debatten .
Jag förklarar debatten för avslutad .
Omröstningen kommer att äga rum nu .
Förslag till gemensam resolution om skydd för biståndsarbetare .
( Parlamentet antog resolutionen . )
Röstförklaringar Herr talman !
Jag avstod från att rösta eftersom jag anser att det är nödvändigt att man från kommissionens sida fortsätter sina intensiva kontakter med regeringen , men å andra sidan också anstränger sig för att arbeta intensivare tillsammans med de icke-statliga organisationerna .
Jag tror att mediapolitik också är mycket viktig , att vi också informerar befolkningen på platsen om vad som faktiskt sker .
Det bör även vara vår politik att föra samman de båda stridande parterna .
Här har kommissionen redan gjort väldigt mycket , och jag önskar den för detta allt gott för framtiden !
Herr talman !
Jag röstade för detta förslag om skydd för biståndsarbetarna i världen eftersom jag anser att det är en viktig uppgift för Europeiska gemenskapen att försvara de egna biståndsarbetarna som över hela världen utför ett så viktigt arbete .
Europeiska unionen borde skapa regler på detta område .
Jag hoppas att kommissionen inser att när man bedriver handel med alla stater så måste man också begära att frivilligarbetarna får hjälp och skydd och man måste agera så att den som reser för att hjälpa medborgare i andra länder är väl förberedd , utbildad och skyddad och att vederbörande ges en möjlighet att fullfölja sin uppgift .
Europeiska unionen får inte glömma bort dem bland de egna medborgarna som utför ett så viktigt arbete över hela världen .
Ärade kollegor , alla punkter på dagordningen är genomgångna .
Protokollet från sammanträdet kommer att underställas parlamentet för godkännande i början av nästa sammanträdesperiod .
 
Avbrytande av sessionen Jag förklarar Europaparlamentets session avbruten .
( Sammanträdet avslutades kl .
10.40 . )
