 
Justering av protokollet från föregående sammanträde Protokollet från föregående sammanträde har delats ut .
Finns det några synpunkter ?
Herr talman !
Jag svarar på en uppmaning från parlamentets talman i går eftermiddag att för min grupps räkning tala om ett ärende som det hänvisas till i protokollet .
Jag syftar på punkt 11 på föredragningslistan .
För det första , anser jag att den fråga som socialistgruppens ordförande tog upp i går om att återinsätta debatten med kommissionens ordförande om det femåriga strategiska programmet var tillräckligt viktig för att andra talare som kort ville kommentera denna fråga skulle kunna tillmötesgås .
Jag vill uttrycka denna uppfattning även om jag med all respekt inte instämde i utan röstade emot socialistgruppens ordförandes förslag .
Det andra påpekande jag skulle vilja göra - och som jag skulle ha velat göra i går före omröstningen - är att detta parlament som andra talare kommenterade i går bara kan åstadkomma någonting genom ett nära samarbete med Europeiska kommissionen som ger synergieffekter .
Vi bör också vara ödmjuka nog att erkänna att vi , om vi hade velat ha en strategisk debatt som inte bara åtföljdes av en föredragning och ett klargörande av kommissionens ordförande utan också av ett femårsprogram , skulle ha haft strukturerna på plats långt tidigare än en vecka innan debatten i denna kammare , så att vi hade kunnat diskutera och i sinom tid meddela kommissionen våra önskemål .
Det finns en grundläggande lärdom jag skulle vilja att vi drog av detta .
När större viktiga debatter är inplanerade mellan denna kammare och Europeiska kommissionen i framtiden bör vi reda ut vilka våra ömsesidiga förväntningar är , åtminstone en hel arbetsmånad i förväg .
Först och främst krävs klarhet mellan alla grupper i denna kammare och sedan mellan detta parlament och kommissionen .
Vi bör inte för sent upptäcka att vi befinner oss i den olyckliga positionen att en eller annan institution skapar en onödig spricka i relationerna mellan institutionerna .
När man läser några av pressens rapporter från i fredags verkar det som om kommissionen och dess ordförande utövade en lovvärd självkontroll i sina offentliga kommentarer .
Detta är någonting jag uppskattar mycket .
Jag hoppas att vi kommer att lära oss läxorna och inte upprepa denna onödiga övning , som jag tror berodde på ett missförstånd om vad som förväntades och inte på ond tro hos någon av de två institutionerna .
Det bör inte förstoras till någonting mer än så .
( Applåder ) Tack så mycket , herr Cox !
Jag förstår vad ni menar .
Vi har noterat det .
Herr talman !
Beträffande punkt 11 i arbetsplanen kom vi i går överens om att Bourlanges betänkande skulle vara med på dagens föredragningslista .
Emellertid drogs det tillbaka av budgetutskottet i går kväll utan att diskuteras eller bli föremål för omröstning .
Det måste därför strykas från dagens föredragningslista . .
Herr Wynn , det är logiskt .
Betänkandet har följaktligen avförts från föredragningslistan .
Herr talman !
Vad beträffar Lynnes kommentarer i går om hälsa och säkerhet i denna byggnad antar jag att hon talade om avloppet , för det finns en hemsk kloaklukt på femte våningen i tornet .
Detta måste undersökas eftersom det är ett klart tecken på att någonting är väldigt fel .
Jag vill inte komma dragande med frågan om denna byggnad i all oändlighet , men detta är ett allvarligt problem . .
Fru Ahern , vi har noterat det .
Jag vill be er att lägga fram detta speciella fall , som rör fläktarna på en viss våning , för kvestorerna , eftersom de egentligen är ansvariga för det .
Men vi skall också vidarebefordra det till våra enheter .
Tack så mycket !
( Parlamentet justerade protokollet . )
 
Reformering av den europeiska konkurrenspolitiken Nästa punkt på föredragningslistan är gemensam debatt om följande betänkanden : A5-0069 / 1999 av von Wogau för utskottet för ekonomi och valutafrågor om kommissionens vitbok om modernisering av reglerna om tillämpning av artiklarna 85 och 86 i EG-fördraget ( KOM ( 1999 ) 101 - C5-0105 / 1999 - 1999 / 2108 ( COS ) ) , A5-0078 / 1999 av Rapkay för utskottet för ekonomi och valutafrågor om den XXVII : e rapporten om konkurrenspolitiken ( 1998 ) ( SEK ( 1999 ) 743 - C5-0121 / 1999 - 1999 / 2124 ( COS ) ) , A5-0087 / 1999 av Jonckheer för utskottet för ekonomi och valutafrågor om sjunde översikten över statligt stöd i Europeiska unionen inom tillverkningsindustrin och vissa andra sektorer ( KOM ( 1999 ) 148 - C5-0107 / 1999 - 1999 / 2110 ( COS ) ) , ( rapport 1995-1997 ) , A5-0073 / 1999 av Langen för utskottet för ekonomi och valutafrågor om kommissionens rapport om 1998 års genomförande av kommissionens beslut nr 2496 / 96 / EKSG av den 18 december 1996 om gemenskapsregler för statligt stöd till stålindustrin ( gemenskapsreglerna för stöd till stålindustrin ) ( KOM ( 1999 ) 94 - C5-0104 / 1999 - 1999 / 2107 ( COS ) ) . .
( DE ) Herr talman , mina damer och herrar , kära kolleger !
Kommissionens vitbok om modernisering av de europeiska konkurrensreglerna har utlöst en intensiv och livlig debatt bland den intresserade allmänheten .
Reaktionerna från experter och berörda parter sträcker sig från totalt avvisande till förbehållslöst stöd .
Vad handlar det nu om i denna vitbok ?
Det befintliga systemet med de europeiska konkurrensreglerna inrättades under gemenskapens första år .
Detta system , som är baserat på ett centraliserat anmälnings- och godkännandeförfarande , var säkert bra under de villkor som då rådde .
Detta förfarande har väsentligt bidragit till att skapa en europeisk konkurrenskultur .
Under de 40 år som gått sedan det skapades har emellertid ramvillkoren väsentligt förändrats .
De sex länderna i gemenskapen har utökats till 15 , och står inför en ytterligare utvidgning till 27 medlemmar .
Systemet är dock till största delen likadant .
Det är därför absolut nödvändigt med en reform .
Detta bestrids heller inte från något håll i debatten .
Visserligen anser vissa kritiker att kommissionen går alltför långt med sina förslag .
Kommissionen vill avskaffa systemet med anmälningar och godkännanden , och i stället stärka de nationella myndigheternas och domstolarnas roll vid tillämpningen av konkurrensreglerna .
Det handlar med andra ord om övergång från ett godkännandesystem till ett system med direkt tillämplighet av undantagsregeln .
Förbudsprincipen - och detta är viktigt - bibehålls dock .
Principiellt anser jag att om en myndighet som påstås ha en tendens till byråkrati och centralism kommer med ett förslag om en avbyråkratisering och en decentralisering bör vi åtminstone allvarligt granska detta förslag .
Enligt kommissionens förslag handlar det enbart om de konkurrensbegränsande överenskommelserna mellan företag liksom om missbruk av dominerande ställning .
Anmälningsplikten vid statligt stöd och företagssammanslutningar bibehålls dock .
Utskottet för ekonomi och valutafrågor har principiellt godkänt dessa förslag från kommissionen med endast en röst emot och två nedlagda röster .
En avslutande bedömning kommer dock att vara möjlig först när kommissionen lägger fram de lagförslag som nu förväntas .
Även om jag principiellt röstar för kommissionens förslag , finns det dock en rad punkter som behöver förbättras eller åtminstone klargöras .
Några av dessa punkter vill jag kortfattat förklara .
Flera kritiker av vitboken menar att decentraliseringen äventyrar samstämmigheten i gemenskapens rättstillämpning .
Nationella myndigheter och i synnerhet domstolarna skulle ännu inte överallt vara i stånd att spela den roll som kommissionen avser när det gäller att tillämpa konkurrensreglerna .
För det första har de nationella kartellmyndigheterna under det senaste årtiondet blivit tillräckligt förtrogna med tillämpningen av konkurrensreglerna .
För det andra har de nationella domstolarna redan i enlighet med nuvarande rättsskipning behörighet att tillämpa artiklarna 81.1 , 82 och 86 .
Trots detta är det fortfarande mycket viktigt att kommissionen stöder de nationella myndigheterna och domstolarna med gruppundantagsförordningar , riktlinjer och meddelanden .
Dessutom måste samarbetet mellan de nationella myndigheterna och kommissionen stärkas , liksom mellan de nationella myndigheterna .
Vad beträffar de nationella domstolarnas behörighet föreslår vi i föreliggande betänkande att det föreskrivs domstolar som är specialiserade på konkurrensrättsligt förfarande .
Detta praktiseras redan nu med framgång i vissa medlemsländer .
Från företagarnas sida befaras att man skall förlora i rättssäkerhet .
För att motverka detta bör företagen i vissa fall få behålla möjligheten att erhålla ett förhandsgodkännande från kommissionen .
Detta är endast några , ehuru centrala aspekter , som man måste ta hänsyn till vid moderniseringen av de europeiska konkurrensreglerna .
Vi befinner oss fortfarande bara i början av förfarandet .
Diskussionen kommer att fortsätta tills man slutligen kommer fram till konkreta lagförslag .
Med vitboken är vi dock - det är jag övertygad om - på rätt väg .
Under de gångna årtiondena har en europeisk konkurrenskultur utvecklats .
Den av kommissionen föreslagna decentraliseringen svarar mot subsidiaritetsprincipen , som ju nu också är förankrad i fördraget .
Detta leder till en ökad tillämpning av de europeiska konkurrensreglerna på nationell och regional nivå och gör det möjligt att bredda grundvalen för den europeiska konkurrenskulturen .
Avslutningsvis vill jag säga att den reformering av konkurrenspolitiken , som här inleds , är nödvändig , och att det är särskilt nödvändigt att klargöra att Europeiska unionens konkurrenspolitik är en väsentlig förutsättning för att man skall lyckas med en marknadsekonomi med socialt ansvar .
Både kommissionen och parlamentet måste på ett tydligare sätt än hittills klargöra att konkurrenspolitiken , konkurrensen mellan företagen och det faktum att kommissionen vakar över den , hör till det medborgarna är främst intresserade av .
( Applåder ) Herr talman , herr kommissionär !
Vi för i dag en viktig debatt om Europeiska unionens konkurrenspolitik .
Vi diskuterar en mycket omstridd modernisering av den europeiska kartellrätten , nämligen Wogaus betänkande , och den är mycket mer omstridd än kanske omröstningen i utskottet för ekonomi och valutafrågor gett vid handen .
Jag vill absolut säga att jag personligen anser att kommissionens förslag i detta konkreta fall är felaktigt , och att det återstår att se huruvida begreppet modernisering verkligen är befogat för vitbokens innehåll i artiklarna 81 och 82 , eller om inte snarare begreppet tillbakagång vore mer tillämpligt i detta fall .
Vi talar i dag emellertid också om översikten över statligt stöd och den allmänna rapporten om konkurrenspolitiken för 1998 , där mitt inlägg i denna gemensamma debatt gäller det senare området .
Men båda områdena - rapporten om konkurrenspolitiken och översikten över det statliga stödet - har naturligtvis också en gemensam grundval i denna vitbok .
Det gäller kravet på modernisering , på den europeiska konkurrenspolitikens framtidsförmåga .
Om man läser kommissionens båda dokument ser man att 1998 var ett år där man fortsatt den modernisering som inletts under 1997 och delvis också avslutat den ; det känner vi själva till från vårt löpande parlamentariska arbete .
Låt mig göra två principiella påpekanden : Kommissionen har , som ansvarig myndighet , med sin konsekventa hållning alltid gjort stora insatser för konkurrensfriheten , inte alltid till glädje för berörda medlemsstater eller företag .
Den bör fortsätta på denna väg .
Men , herr kommissionär , allt detta blir i framtiden inte mindre komplicerat - jag vill bara erinra om utmaningarna på grund av utvidgningen av unionen , fördjupningen av den inre marknaden , de tekniska framstegen och globaliseringen .
Det hänger faktiskt inte bara på moderniseringen av gemenskapsrätten , utan det beror mer än någonsin på öppenheten i besluten i de enskilda fallen , och på möjligheten att även kunna sätta sig in i besluten , ty den europeiska konkurrenspolitiken kommer att vara beroende av acceptansen från befolkningen , liksom från de berörda politiska instanserna och företagen .
Men - utan öppenhet ingen acceptans , och då alltså inte heller någon modernisering utan öppenhet .
Rapporten om konkurrenspolitiken 1998 är inte någon dålig grundval för detta , men det finns inte heller någonting som inte skulle kunna göras bättre .
En rad impulser kommer vi att lämna vidare till er , herr kommissionär , tillsammans med vår resolution , men en delaspekt vill jag redan nu gå in på : Öppenhet och redovisningsskyldighet hör ihop .
Jag vill inte rubba ansvarsfördelningen mellan kommissionen och parlamentet .
Kommissionen är det verkställande organet , och parlamentet bör för sitt eget oberoendes skull inte heller vilja vara det , utan parlamentet är ett kontrollorgan , och var kan man bättre klargöra bakgrunden till sina beslut än i det demokratiskt valda parlamentet och just i en ständig parlamentarisk diskussion ?
Även här bör vi fortsätta på den inslagna vägen , intensifiera den och göra den beständig .
Men en sak vill jag säga helt tydligt : Parlamentet är lagstiftande , och att vi just när det gäller konkurrensrätten bara har samrådsrättigheter , är egentligen skandal !
Här riktar vi ett krav till rådet och regeringskonferensen att införa ett medbeslutandeförfarande när det gäller konkurrensrätten .
Jag förväntar mig av kommissionen att man fullständigt utnyttjar alla möjligheter till parlamentarisk medverkan , om det finns tvivel om att parlamentet skall kunna delta , och detta också redan i den fördragssituation vi har nu .
Jag förväntar mig också att kommissionen kommer att stödja oss offensivt i fråga om kravet på medbeslutande i lagstiftningsförfarandet .
Det kommer att utgöra ett prov på hur klokt våra institutioner kan samarbeta .
Trots att man bekänner sig till konkurrensprincipen är konkurrensen dock inte något mål i sig .
Konkurrens är ett instrument och leder inte alltid till optimala lösningar .
Det hör nu en gång till de elementära kunskaperna i ekonomi att marknaden i många avseenden misslyckas , och den som bestrider detta är en ideolog , och ingenting annat .
Konkurrensen skall balansera utbud och efterfrågan , och sörja för en optimal fördelning av de ekonomiska resurserna .
Men en optimal effektivitet inställer sig inte nödvändigtvis av sig själv .
Det krävs ramvillkor för att förhindra missbruk , till exempelvis genom kartellrätten .
Men därmed förhindras huvudsakligen endast missbruk , det räcker inte ensamt till för att uppnå de mål som legitimeras av samhället .
Ja till konkurrens , och en inskränkning av stöden där så krävs och där det är möjligt !
Men eftersom stöden i rapporten om konkurrenspolitiken 1998 utgör den största delen vill jag , oaktat kollegan Junkers betänkande , ändå tillfoga följande : Stöd till små och medelstora företag när det gäller forskning och utveckling , när det gäller utbildning i regionalpolitik och miljöpolitik , det är absolut möjligt och måste också vara genomförbart .
Stöd måste tillåtas just för sådana mål , så länge de inte leder till oacceptabla snedvridningar av konkurrensen .
Just här är det ännu viktigare att besluten är förståeliga än i fråga om kartell- och fusionsrätten .
Stöden bör inte nedvärderas , utan man måste se på hur de kan bidra till att man uppnår de mål som just nämnts .
Det sista påpekandet riktade sig mindre till kommissionen , utan snarare till kollegerna i PPE-gruppen .
Herr talman , herr kommissionär , mina kära kolleger !
Det betänkande som jag i dag har tillfälle att lägga fram för er , är ett yttrande om kommissionens årliga rapport över statliga stöd inom Europeiska unionen , för vilka gemenskapen är behörig i kraft av artiklarna 87 , 88 och 89 i fördragen .
Kommissionens rapport är i huvudsak beskrivande ; här redogörs för statsstödens utveckling såväl inom tillverkningsindustrin som inom andra sektorer , enligt kriterier som finansieringsmetoder och eftersträvade mål .
När det gäller rapportens kvantitativa avsnitt tillåter jag mig att hänvisa till motiveringen .
Här nöjer jag mig med att peka på att årsbeloppet i genomsnitt ligger på 95 miljarder euro för perioden i fråga , vilket utgör en minskning på 13 procent i förhållande till perioden 1993-1995 , något som i huvudsak beror på en minskning av stöden i Förbundsrepubliken Tyskland .
I klartext ligger de anmälda statsstöden i stort sett på ett stabilt genomsnitt under den granskade perioden , och tar ungefär 1,2 procent av gemenskapens BNI i anspråk .
Det motsvarar händelsevis mer eller mindre gemenskapens budget för ett år .
Samtidigt är skillnaderna mellan staterna avsevärda och kan bedömas på olika sätt , bl.a. i procent av mervärdet och per löntagare .
Det kan också vara av intresse att lägga till de statliga stöd och gemenskapens interventioner som på något sätt kan likställas med statsstöd .
Då framgår det klart och tydligt att det är de fyra länder som bl.a. får stöd från Sammanhållningsfonden som hamnar i toppen av klassificeringen .
Därmed kommer jag fram till betänkandets förslagsdel .
Vi kan först och främst konstatera att kommissionen anser att informationen ( såsom den presenteras i kommissionens årliga rapport ) täcker alltför stora områden för att tillåta en grundligare utvärdering av statsstödspolitiken , något som är såväl berättigat som förnuftigt med hänsyn till nationella intressen , och mycket viktigt med avseende på respekten för konkurrensen , enligt definitionen i fördragets bestämmelser .
Kommissionen kan endast samla in och analysera de uppgifter som medlemsstaterna anmäler .
Det är således staternas och regionernas sak att garantera kvaliteten på de uppgifter som lämnas in , och vårt utskott anser att man bör göra ytterligare insatser för det ändamålet .
Av samma skäl försvarar vårt parlamentsutskott det redan gamla förslaget om ett offentligt register över statsstöden , som bl.a. skall finnas tillgängligt på Internet .
Om uppgifterna blir bättre och mer detaljerade , i synnerhet i förhållande till eftersträvade mål och noterade resultat , kommer Europeiska kommissionen själv att kunna företa , eller låta företa , regelbundna studier för en social och ekonomisk utvärdering av nationella och regionala stöd .
I den mån sådana studier redan finns , bör kommissionen så öppet som möjligt informera om dess egna synpunkter i förhållande till fördragens mål , som inte bara är att säkerställa den europeiska ekonomins konkurrenskraft , utan också en hållbar utveckling och ekonomisk och social sammanhållning .
Genom att i första hand lägga tonvikt på kvaliteten på den information som lämnas , har vårt utskott undvikit att - i våra debatter och därmed i det betänkande som jag har äran att presentera för er - göra det enkelt för oss genom att i förväg hävda att statsstöden i sig är alltför stora alternativt otillräckliga .
En majoritet av utskottets ledamöter har i stället strävat efter en jämvikt ; å ena sidan bör man kräva att såväl staterna som företagen respekterar konkurrensreglerna och å andra sidan bör man erkänna att den här typen av stöd kan medverka till att fördragets mål förverkligas , i synnerhet , som jag redan har nämnt , i fråga om hållbar utveckling , forskning och utveckling samt ekonomisk och social sammanhållning .
Samtidigt har utskottet godkänt en rad olika ändringsförslag till föredragandens ursprungliga utkast , vilka bl.a. betonar att stöd som bedöms vara illegala skall betalas tillbaka och att det upprättas en resultatlista .
Sju ändringsförslag har givits in på nytt inför det här plenarsammanträdet .
Flertalet av dem förmedlar våra politiska skiljelinjer i fråga om statsstödens lämplighet och effektivitet , med tanke på att enbart privata investeringar inte räcker till , vare sig detta medges eller ej , market failures eller marknadens otillräcklighet .
Det finns bl.a. ett ändringsförslag rörande energisektorn , som jag i egenskap av föredragande vill framhålla som särskilt betydelsefullt .
Herr kommissionär !
Jag vill avsluta denna presentation genom att å ena sidan framhålla ett orosmoln och å andra sidan en begäran från ledamöterna i vårt utskott .
Oron avser de central- och östeuropeiska ländernas anslutningsprocess i förhållande till konkurrenspolitik och statsstöd .
Detta är med största sannolikhet en komplicerad fråga , och vi skulle önska att kommissionen redogjorde för sakens nuvarande läge , bl.a. vad gäller de ansökande ekonomiernas kapacitet att respektera konkurrensreglerna , och när det gäller statsstöd ; det sannolika behovet av att fastställa specifika regler om statsstöd för en omstrukturering av deras sektorer .
Till sist , och härmed skall jag avsluta , en begäran som rör Europaparlamentets framtida behörighet inom de områden som vi nu talar om - konkurrenspolitik och statsstöd - en möjlighet med tanke på nästa regeringskonferens .
Som ni vet , herr kommissionär , försvarar vi i detta betänkande tanken att medbeslutandeförfarandet skall tillämpas för grundläggande lagstiftning om statliga stöd . .
( DE ) Herr talman , herr kommissionär , mina damer och herrar !
Min del i dagens debatt gäller gemenskapsreglerna för stöd till stålindustrin .
Det är det allmänna stödet som lämnats i Europa i enlighet med dessa gemenskapsregler , och som kommissionen har granskat .
Det är totalt 27 fall under år 1998 .
Dessa fall har kommissionen avgett en egen rapport om .
EKSG-fördraget kommer att löpa ut inom kort .
Den fråga som vi i dag i synnerhet måste ägna oss åt är hur stödet till stålindustrin skall hanteras i framtiden .
Kommissionens beslut , som framläggs i översikten , välkomnas av Europaparlamentet , inklusive beslutet att i ett konkret fall kräva tillbaka medlen med tillämpning av artikel 88 i EKSG-fördraget .
Den europeiska stålindustrins konkurrenskraft behandlas samtidigt också i kommissionens senaste meddelande , som vi ännu inte har diskuterat i parlamentet .
Liksom på andra områden gäller även för järn- och stålindustrin ett generellt förbud mot stöd enligt artikel 87.1 i EG-fördraget .
Enligt denna artikel är statligt stöd principiellt oförenligt med den gemensamma marknaden .
Undantag tillåts endast i exakt definierade fall .
Enligt artikel 88 är kommissionen ålagd att kontrollera statliga stöd .
År 1998 var det viktigaste fallet när Preussag i Tyskland försågs med kapital till ett belopp av 540 miljoner euro .
Dessutom måste medlemsstaterna meddela kommissionen sina stödåtgärder i förväg .
Vad beträffar stålindustrin ställdes de gällande reglerna upp den 18 december 1996 .
Enligt dessa kan stöd till förmån för stålindustrin endast lämnas i bestämda , exakt definierade fall .
Det är forsknings- och utvecklingsstöd , miljöskyddsstöd , socialt stöd vid stängning av stålverksanläggningar och stöd för den slutliga nedläggningen i icke konkurrenskraftiga företag .
Dessutom finns det en särbestämmelse om upp till 50 miljoner euro för medlemslandet Grekland .
Uppenbarligen har det under de gångna åren ändå uppstått problem i den praktiska hanteringen av gemenskapsreglerna till stöd för stålindustrin , som inte har tagits upp fullständigt i betänkandet .
Ur parlamentets synvinkel är det viktigt att man redan i dag talar om bestämmelser som kan träda i kraft när dessa gemenskapsregler för stöd till stålindustrin har löpt ut .
Det får inte beslutas om någon uppmjukning av befintliga grundvalar för gemenskapsreglerna för stöd till stålindustrin .
Ingen vill ha en hämningslös subventionskonkurrens i Europa .
Detta skulle avsevärt skada den inre marknaden även efter den konsolidering av stålindustrin som skett under de senaste åren .
Därför anser parlamentet att det är nödvändigt att bestämmelserna om subventioner till stålindustrin ändras med tanke på skillnad i behandling som industrin påstår har ägt rum , och att kommissionen för rådet lägger fram bestämmelser som skall träda i kraft när de nuvarande bestämmelserna löpt ut .
Vi känner till att rådet hittills vägrat besluta om sådana bestämmelser .
Det beror också på att man tror att man , när gemenskapens regler om stöd till stålindustrin löper ut , återigen kan göra som man vill , utan den besvärliga kontrollen från kommissionens sida .
Vi kräver därför att gemenskapsreglerna om stöd till stålindustrin skall regleras genom en förordning från rådet enligt artikel 94 när fördraget löpt ut , eftersom de endast på så sätt kan bli klara och rättsligt bindande .
Det strikta förbudet mot allt stöd , som inte täcks av gemenskapsreglerna , kan bara iakttas på detta sätt .
En förordning från rådet , som omedelbart träder i kraft , måste också iakttas av de regionala regeringarna .
Även i framtiden måste vi undvika intrång i konkurrensvillkoren och störningar i balansen på marknaderna .
Man måste också kritisera kommissionens praxis att godkänna upprepat stöd för stålföretag , som enligt kommissionens åsikt inte faller under kategorierna i gemenskapsbestämmelserna , även om EG-domstolen i enstaka beslut har godkänt denna skillnad i behandling .
I ett betänkande som återstår att utforma för år 1999 uppmanas kommissionen att detaljerat klarlägga sin aktiva roll vid utarbetandet av omstruktureringsplaner och godkända undantagsfall , och därmed på denna grundval möjliggöra en korrekt utvärdering av de totala sammanhangen .
Efter att utskottet för ekonomi och valutafrågor enhälligt har antagit förslaget till betänkande , med två nedlagda röster , ber jag att vi i kammaren helt och fullt godkänner denna framställning , som vi själva har initierat . .
Herr talman , kära kolleger !
Den inre marknaden är inte fullbordad .
Subventioner , monopol och konkurrenshinder hämmar fortfarande både marknader och utveckling .
Nationella regeringar skjuter till subventioner och lovar att det är sista gången , men så upprepas det igen .
Subventioner snedvrider allokeringar , både inom och mellan länder .
En successiv avveckling av statsstödet behövs , och alltfler marknader måste öppnas för konkurrens .
Det gäller både dem som har monopoliserats privat och offentligt .
Offentliga monopol avvecklas oftast motvilligt .
Ökad konkurrens och nyetableringar skulle kunna ge betydande välfärdsvinster - även inom utbildning , sjukvård och social service .
Offentliga monopol måste ersättas av konkurrenskraftiga strukturer .
Europa måste moderniseras och anpassas till entreprenörskap och en konkurrenskraftigare miljö för konsumenter och företag .
Effektiv konkurrens pressar priser och höjer levnadsnivåer .
Konsumentpolitiken har i alltför liten utsträckning inriktat sig på just prisnivåerna .
Konkurrenspolitik och konsumentpolitik hör ihop .
Inre marknaden är grunden för vårt arbete .
Dess lagstiftning skall gälla lika för alla , för stora som för små länder .
En systematisk genomgång av de nationella regelverken behövs för att undanröja konkurrenshinder .
Även EU : s eget regelverk kan då behöva en analys .
Den nya modell som nu prövas av kommissionen får inte leda till en ren nationaliseringsprocess som skulle urholka den uppnådda konkurrenspolitiken .
Den måste vara väl förankrad i medlemsstaternas nationella myndigheter för att bli effektiv .
Om ett halvår kan det vara lagom att göra en analys av utfallet , men även att se närmare på den nya situationens effekter på kommissionens roll .
Tanken på att hålla en institutionellt övergripande kongress som öppnar för en förutsättningslös debatt utifrån ett brett perspektiv med representanter från olika intressenter har tills vidare löst frågan om hur man skall gå vidare .
Då finns det tillfälle att slå fast nya principer eller återkomma till de mer genomgripande förändringar som har diskuterats .
Då gives också tillfälle att finna nya gemensamma lösningar och analysera ändringsförslagen från utskottsdebatten .
Rättstillämpningen i konkurrensfrågor måste vara korrekt .
Felaktigt tillämpad konkurrenspolitik kan orsaka rättsförluster och göra ingrepp i äganderätten , vilket är en viktig , grundläggande princip som vi skall slå vakt om .
Det ligger en ganska spännande debatt framför oss .
En konferens där frågorna ventileras möjliggör att missförstånd kan rätas ut , samtidigt som vissa punkter också kanske kan förbättras .
Parlament och kommission kan tillsammans stärka insatserna för en effektiv konkurrenspolitik och därmed skapa nya möjligheter och nya resurser för medborgarna .
Just i min valkrets , Stockholm , har vi många goda lokala exempel på ökat utbud och förbättrad kvalitet som uppstått just på grund av konkurrensutsättningar på tidigare helt monopoliserade områden .
Vi tillskyndar en fortsättning på den öppna debatt som stärkts under behandlingen av betänkandena av von Wogau och Rapkay .
Vi hoppas att de rättsliga synpunkterna också kommer att tillmätas den vikt som är rimlig i en rättsstat .
Herr talman , kära kolleger !
Det gläder mig att jag får hålla mitt första tal här i dag som ny ledamot , även om det sker med en viss försening .
Först vill jag tacka föredragandena von Wogau , Langen , Rapkay , Jonckheer samt kommissionen för det mycket goda samarbetet .
Konkurrensen utgör säkerligen grundvalen för en marknadsekonomi med socialt ansvar , och den europeiska konkurrenspolitiken har varit framgångsrik , inte minst vad gäller energi och telekommunikation , och har lett till märkbart lägre priser och bättre service .
Allt till konsumenternas fördel .
Men nu har vi kommit fram till en punkt där vi måste vidareutveckla konkurrenspolitiken .
Här har kommissionen lagt fram en ny vitbok med två kärnpunkter : Anmälningsplikten skall överges , och den rättsliga verkställigheten skall återföras .
Att man överger anmälningsplikten innebär i varje fall mindre byråkrati och administrativa kostnader .
Denna systemändring leder naturligtvis samtidigt till mer ansvar för de enskilda i näringslivet .
Det är inte längre så enkelt att man bara lägger fram något och får det godkänt , utan nu måste alla till att börja med själva bära ansvaret , och det är kanske också orsaken till att en eller annan där ute uppfattar detta som obehagligt .
Men jag tror att vi bör utnyttja chansen att låta Europa också ge en signal till mindre byråkrati .
Den andra punkten är återföringen av den rättsliga verkställigheten .
För att en rättslig kultur skall kunna skapas i Europa måste rätten givetvis inte bara tillämpas av kommissionen och av centrala organ , utan också av nationella myndigheter och domstolar .
Vi säger ju inte heller att all EG-rätt alltid skall beslutas centralt , men just i anpassningsfasen kommer det att finnas en viss osäkerhet vad gäller rätten .
Här är det säkerligen nödvändigt , i det lagstiftningsförfarande som vi står inför , att utveckla ett instrument för att ge företagen rättssäkerhet och möjlighet att vända sig till kommissionen .
Det bör hållas en dörr öppen till en europeisk kartellmyndighet , som säkert kommer att diskuteras i framtiden .
Men vi behöver mer öppenhet i konkurrenspolitiken .
Parlamentet måste bli mer delaktigt , och jag tror också att om vi inför ett register , där vi kan se vilka statliga åtgärder som vidtas , så kommer detta att leda till disciplinering i medlemsstaterna .
Vad gäller konkurrensen i framtiden ligger emellertid två punkter mig mycket varmt om hjärtat .
Det ena är subsidiariteten .
Vi anser alla att konkurrens är nödvändig för ekonomin och främjar prestationsförmågan , och jag tror att vi också bör släppa in konkurrens i regionerna .
Konkurrensen mellan regionerna kommer säkerligen att stärka Europeiska unionen , och inte försvaga den .
Här kan jag nämna exemplen med GA-stöd , sparkassor och delstatsbanker , samt kvalitetsgaranti .
Här har en region av egen kraft skapat något för att saluföra sina egna produkter .
Dessa egna initiativ får inte förstöras från europeiskt håll .
Jag tror att det också är nödvändigt med en höjning av Deminimus-bestämmelserna .
Vi bör satsa allt på att påskynda konkurrensen mellan regionerna .
Det andra är en diskussion om konkurrens och marknadsekonomi med socialt ansvar , och då talar jag här inte om misslyckanden från marknadens sida .
Jag har ju redan nämnt exemplen med delstatsbanker och sparkassor , men jag vill driva det som man alltid hör från det ena eller andra hållet till sin spets .
En boende på ett ålderdomshem är i dag socialt placerad .
Men man kan också betrakta honom som en kund , och jag tror att vi ganska tydligt och i god tid bör diskutera var det sociala området , var de strukturer som vuxit upp sätter stopp för konkurrensen .
Annars kan jag här använda uttrycket kunder för detta område , och därigenom mycket starkt förstöra sociala områden .
Slutligen vill jag också säga i fråga om subsidiaritetsprincipen : Jag anser att det är absolut nödvändigt att där medlemsländerna medger att regioner och kommuner kan uppbära skatter skall detta bibehållas och inte regleras enhetligt av Europa . .
Tack så mycket , herr kollega .
Jag gratulerar er till det som man inom den tyska parlamentarismen , i ert fall felaktigt , kallar för ett jungfrutal .
Herr talman , herr kommissionär , kära kolleger !
Jag kommer att tala å min kollega Robert Goebbels vägnar , eftersom han inte kunde komma på grund av politiska förpliktelser .
Inom utskottet för ekonomi och valutafrågor väckte Jonckheerbetänkandet bittra kontroverser kring marknadens sätt att fungera .
En knapp högermajoritet lyckades stryka samtliga hänvisningar till att marknaden har brister .
Men även om majoriteten i vårt parlament skulle följa denna ultraliberala uppfattning om en så kallad perfekt marknad , skulle världen inte förändras för det .
Ekonomiska rapporter från den verkliga världen ger tillräckliga bevis för att man inte på något sätt skapar en perfekt konkurrens och bästa möjliga resursfördelning genom att avskaffa alla former av offentliga interventioner på marknaden .
Marknaden må ha varit människors främsta handelsplats sedan urminnes tider , men den har aldrig varit perfekt .
Marknaden gynnar kortsiktighet och omedelbara vinster .
På marknaden verkar styrkeförhållandena mellan utbud och efterfrågan i allmänhet till de svagares nackdel , konsumenterna , arbetarna .
För att fungera fordrar marknaden regler .
Den nödvändiga och värdefulla initiativandan måste åtföljas av en känsla av ansvar gentemot samhället .
Vi europeiska socialister är för en marknadsekonomi med sociala ändamål .
Marknaden är inte ett mål i sig ; den skall bidra till att förbättra de mänskliga villkoren .
Europeiska unionen och staterna skall inte ta de ekonomiska aktörernas plats , men statsmakterna måste fastställa regler och mål som gör att ekonomin kan utvecklas på ett hållbart sätt .
Statliga stöd kan slutligen möjliggöra omstruktureringar , erbjuda utbildning , rädda arbetstillfällen och därmed kunnande .
Huvudmålet med unionens konkurrenspolitik får inte vara att minska den allmänna stödnivån .
De statliga stöden måste anpassas efter unionens mål , framför allt ekonomisk och social sammanhållning , hållbar utveckling samt forskning .
Kommissionen måste bedriva klappjakt på illegala stöd och de stöd som verkligen blockerar den inre marknaden .
Men att avskaffa alla former av statsstöd skulle vara ett allvarligt misstag .
Internet är inte en marknadsprodukt , utan resultatet av forskning som finansierats av den amerikanska armén .
World Wide Web , som har möjliggjort en blixtrande utveckling av informationssamhället , utvecklades av Europeiska atomforskningscentret ( CERN ) i Genève , återigen med hjälp av statsstöd .
Att den tyska regeringen räddade Holzmann-gruppen kritiserades som ett ogrundat hinder mot marknadsekonomin .
Centralbankschefen Duisenberg försökte till och med skylla eurons svaghet gentemot dollarn - för övrigt tämligen relativ - på denna statliga interventionism .
Jag har inte hört Duisenberg kritisera det faktum att de amerikanska penningpolitiska myndigheterna räddade Hedge Fund LTCM .
Att vilja rädda 60 000 arbetstillfällen , det är uppenbarligen att begå en synd gentemot marknaden , men att rädda kapital tycks inte skapa några problem för den fria marknadens förespråkare .
Man uppbringar offentliga medel för att reparera de skador som har orsakats av den internationella spekulationen , bl.a. i Mexiko , Asien och Brasilien .
Människors arbete betraktas däremot som vilken justeringsfaktor som helst .
Vi socialister avvisar denna liberala världsfrånvända inställning .
Vi vill ha en riktig konkurrenskultur i Europa .
Den statliga handen måste förbli synlig för att styra marknaden , och kommissionen bör vara dess domare .
Herr talman , bästa kommissionär och kära kolleger !
Jag vill börja med att tacka herr Rapkay för ett väl utarbetat betänkande och ett gott samarbete .
Kommissionär Monti !
Jag vill tacka er för ett utmärkt samarbete och jag vill säga till er att ni nu vid årtusendeskiftet har en mycket viktig funktion .
Ni skall ju städa upp efter de nationella regeringar som har stora visioner på konkurrenspolitikens område , men endast fantasin sätter gränser för vilka olyckor de nationella regeringarna kan åstadkomma .
Jag kan här nämna de senaste exemplen vi har sett : Holzmann , ett företag som fått ett omfattande stöd från den tyska regeringen , sågverk i f.d.
Östtyskland och inte minst stöden till skeppsvarven .
Detta är tre områden inom vilka många danska företag har stora problem och blir utkonkurrerade från marknaden .
Jag vill säga till herr Poos att jag är helt överens med ordförande Duisenberg om att det finns exempel på att några av Europeiska unionens medlemsstater inte är förmögna att omstrukturera sina ekonomier , och därmed bidrar till att undergräva eurons värde .
Den liberala gruppen har lagt fram 80 ändringsförslag i utskottet , som alla rör statligt stöd .
Det är förslag som vi anser leder fram till genomblickbarhet och öppenhet , vilket är mycket viktigt när det gäller att få den inre marknaden att fungera .
Jag vill gärna ta tillfället i akt och tacka mina kolleger i utskottet för deras stöd till den liberala gruppens förslag .
Våra förslag rör som sagt möjligheten till insyn , och jag vill gärna betona det ändringsförslag som uppmanar kommissionen till att utarbeta enhetliga kriterier och villkor för den typ av statligt stöd som vi anser vara lagligt , just för att se till så att företagen kan planera sin situation .
En annan sak är frågan om vad vi skall göra om det statliga stödet förklaras olagligt .
Hur ser vi till att få det olagligt utbetalade statliga stödet tillbaka ?
I dag finns inga gemensamma bestämmelser på detta område och vi uppmanar kraftfullt kommissionen att skapa en harmonisering av bestämmelserna om återbetalning .
Detta är enda sättet för att säkerställa enhetliga konkurrensvillkor .
Till sist föreslår vi att vi dels skapar ett register , vilket flera av mina kolleger varit inne på , men också en resultattavla som visar var länderna står i dag vad gäller statligt stöd .
Ni har visat oss vägen , herr Monti , med en resultattavla för den inre marknaden .
Det är detta som inspirerat oss till att föreslå samma sak vad gäller statligt stöd .
Jag hoppas verkligen att kommissionär Monti kommer att stödja dessa förslag , och jag ser fram emot era kommentarer och er ståndpunkt .
Avslutningsvis vill jag hälsa kommissionens XXVIII : e rapport om konkurrenspolitiken välkommen ; ännu en gång får vi ta del av ett väl utfört arbete .
Men som jag redan har nämnt bör det övergripande syftet fortfarande vara genomblickbarhet och öppenhet .
Det finns fortfarande behov av en uppryckning inom de nämnda områdena och det finns därför en god anledning till att fortsätta med att arbeta på ett målinriktat sätt för att lösa problemen rörande den bristande genomblickbarheten och öppenheten på området för statligt stöd .
Det är inte minst nödvändigt i förhållande till den kommande utvidgningen , och jag vill gärna tacka herr Jonckheer som i sitt betänkande mycket grundligt behandlar problemen i samband med utvidgningen och hur vi skall se till att dessa länder uppfyller våra krav , men också hur vi säkerställer lika konkurrensvillkor .
Det är klar att vi som liberala och gröna har olika uppfattningar om hur vi vill att världen skall se ut , men vad gäller vår målsättning är vi i stort sett överens , och vi vill försöka hitta en förnuftig lösning på våra problem .
Herr talman , herr kommissionär !
Vi har egentligen endast två frågor att svara på .
Är statliga företagsstöd och avtal mellan företag legitima i en marknadsekonomi ?
Och : Vem skall kontrollera undantagen till marknadsekonomins absoluta regler ?
På den första punkten vill vi mycket klart och tydligt säga att det i vissa fall krävs statliga företagsstöd , om vi skall ta hänsyn till de krav på en hållbar utveckling som Europeiska unionen skriver under på , och det oavsett om det sker i form av skattelättnader , differentierad beskattning eller helt enkelt direkta stöd .
Det är också berättigat att det skall kunna finnas avtal och begränsningsavtal mellan företag , eftersom alla sådana avtal bidrar till att dämpa konkurrensens negativa bieffekter på det sociala och miljömässiga planet .
Vi svarar alltså mycket klart och tydligt ja - statliga stöd och avtal är legitima , men vi menar också att varje avtal verkligen måste åtföljas av en motivering .
I von Wogaubetänkandet föreslår man att kontrollen av legitimiteten skall återföras till nationell nivå .
För oss förefaller det ganska riskfyllt , men vi kommer ändå att rösta för , eftersom vi medger att kommissionen inte kan göra allt .
Vi kräver största möjliga öppenhet och att kommissionen skall anförtros största möjliga undersökningsmakt för att i efterhand kontrollera om beviljade undantag är legitima .
Herr talman !
Ännu en gång diskuterar vi Europeiska unionens konkurrenspolitik .
Men under vilka förhållanden förs denna debatt , och vilka slutsatser bör vi komma fram till ?
Dagens verklighet kännetecknas av gigantiska fusioner och sammanslagningar av enorma monopolföretag och skapandet av världsomspännande koncerner med fruktansvärd makt .
Borde vi inte ta upp detta i vår debatt ?
Vilken konkurrenspolitik vill och kan införa kontroller av dessa monopolföretags verksamhet ?
Vissa branscher inom den europeiska industrin , t.ex. varvsindustrin , flygtransporterna , stålindustrin , har drabbats enormt hårt av den konkurrenspolitik som bedrivs .
De har förlorat viktiga marknadsandelar inom världshandeln och hundratusentals arbetstillfällen .
Skall vi inte ta upp detta till diskussion ?
Den skandalösa maktkoncentrationen inom strategiskt viktiga sektorer gör att vinstinriktade multinationella företagsgrupper får kontroll över ekonomin i hela länder - även i unionens medlemsländer .
Trots detta envisas vi med en fortsatt försvagning av den offentliga sektorn , och vi är beredda att skärpa konkurrenspolitiken ytterligare , när vi anser att statliga beställningar från företag av offentlig karaktär också är ett slags statligt stöd .
Å andra sidan leder bortfallet av hundratusentals arbetstillfällen till en våldsam ökning av arbetslösheten .
Arbetstagarna utsätts för ett enormt angrepp på sina arbetsrättsliga och sociala rättigheter .
Konsumenterna ser hur deras levnadsstandard sjunker , hur fattigdomen breder ut sig och hur den offentliga sektorn och den produktiva basen i de flesta av unionens länder skärs ned och upplöses till förmån för en ohämmad och fördärvbringande konkurrens , den totala marknadsekonomin och storkapitalets monopolintressen .
Jag anser att det även är den förda konkurrenspolitiken som bär ansvaret för allt detta , och jag tar fullständigt avstånd från den .
Herr talman , herr kommissionär !
Under brytningsåret , före övergången till den gemensamma valutan , gjorde kommissionen stora ansträngningar för att euron skulle kunna införas under gynnsamma omständigheter .
Konkurrenspolitiken bidrog till denna tilldragelse , inom ramen för dessa medel .
Vi är för vår del fortfarande bestämda motståndare till den gemensamma valutan , som långt ifrån ger oss fördelarna och flexibiliteten med en gemensam valuta , utan i stället stänger in oss i en artificiell tvångsstruktur som påtvingats Europas folk .
Men att styra är samtidigt att förutse och även att ta ansvar , och i det nya framtvingade sammanhanget spelar konkurrensrätten naturligtvis en viktig roll .
På det området har kommissionen prioriterat flera handlingslinjer : att påverka marknadernas struktur genom att aktivt motverka konkurrenshämmande metoder , att inrikta kontrollverksamheten på de affärer som har ett uppenbart gemenskapsintresse samt att markera sin önskan om en modernisering av konkurrensrätten .
Vad gäller statliga stöd måste man se till att bestämmelserna inte blir för tungrodda .
Enligt vår uppfattning är det därför inte önskvärt att införa ett offentligt register över samtliga stöd , eftersom denna tyngande förpliktelse givetvis skulle gå på tvärs mot försöken att lätta på de byråkratiska kraven .
När det slutligen gäller en modernisering av tillämpningen av artiklarna 85 och 86 i fördraget , anser vi inte att en decentraliserad tillämpning nödvändigtvis är ett steg i rätt riktning .
Kommissionen skulle inte endast behålla sin makt att undanhålla de nationella myndigheterna ett ärende - de nationella domstolarna har också klara förpliktelser att undvika varje form av konflikt med kommissionens beslut .
Nationalstaterna skulle således bli kommissionens världsliga rättvisa , med uppdraget att garantera en respekt för tillämpningen av regler som de inte har någon kontroll över .
Sammanfattningsvis vill jag säga att även om vissa bestämmelser går i rätt riktning , kommer vi självklart att förbli vaksamma för att förhindra en federalistisk utveckling , vilket skulle skada Europa och staternas suveränitet .
Herr talman , herr kommissionär , ärade kolleger !
Vi är i allt väsentligt positiva till kommissionens vitbok om konkurrensen , framför allt när det gäller avskaffandet av systemet med meddelande och tillstånd , men vi är också en aning frågande inför ett par punkter .
Framför allt finns risken att delegering av behörigheter till de enskilda staterna , något som i flera avseenden är nödvändigt , kan leda till en alltför kraftig expansion av konkurrensinitiativen och att någon kan frestas att använda antitrustbestämmelserna , inte som en yttersta garanti för att marknaderna skall fungera väl och så som var avsett , utan som ett instrument för den egna ekonomiska och industriella politiken , som ett instrument för planering och ingrepp i marknadernas egna spontana dynamik eller kanske till och med som ett verktyg för protektionistisk politik .
I det avseendet tror jag att vi kan finna vägledning i det som von Eieck har skrivit och säkerligen också i det som den store italienske liberalen Bruno Leoni säger när han just varnar för riskerna för en kraftig ökning av konkurrenshämmande åtgärder .
Det allvarligaste hotet mot marknaden , konkurrensen och valfriheten för de europeiska användarna och konsumenterna är fortfarande hotet om statliga ingrepp i ekonomin .
Det finns statliga stöd till företagen , det har vi redan talat om , det finns fortfarande en stark offentlig närvaro i ekonomin - tänk till exempel på att det italienska finansdepartementet kontrollerar 15 procent av allt kapital på italienska börsen - det finns hinder som regeringar och centralbanker reser inför verksamhet som innebär merger and acquisition ; vi har ofta under de senaste dagarna hört talas om fallet Vodafone-Mannesmann och räddningen av Osman .
Slutligen , herr kommissionär , får vi inte glömma att det fortfarande finns stora ekonomiska sektorer som är i offentliga händer , från den statliga televisionen , som tvångsfinansieras av licensinnehavarna , och postverken , till vissa obligatoriska försäkringssystem , inklusive sjukvårds- och olycksfallsförsäkringar , som hanteras av ineffektiva offentliga monopol som inte ger något val åt användarna om de inte är mycket välbeställda .
Herr kommissionär , jag känner väl till fördragets begränsningar , men jag anser att det även i detta fall är viktigt att understryka att den europeiska ekonomin drabbas hårt av konkurrensen från den amerikanska , även och framför allt på grund av bristen på möjligheter och konkurrens .
Det som vi gör här är förmodligen mycket viktigt , men det är fortfarande otillräckligt .
Herr talman !
Vi för en speciell debatt : om konkurrenspolitik och om statsstöd , statens vänstra och högra hand så att säga .
Medan EMU-kriterierna tvingar medlemsstaterna att begränsa sina utgifter har den höga nivån i fråga om statligt stöd till företagslivet kvarstått .
Förståeligt , för den medlemsstat som börjar med att avveckla statligt stöd löper den största risken att drabbas av företag som flyttar ut , med negativa följder för sysselsättningen .
Men samtidigt obegripligt , för dålig företagaranda och icke livsdugliga arbetsplatser skall inte understödjas med pengar från skattebetalarna .
I princip är enbart horisontala åtgärder tillåtliga eftersom de inte eller knappast rubbar konkurrensen .
Föredragandens ändringsförslag 6 och 7 förtjänar därför stöd .
Ändringsförslagen 1 och 5 visar på fenomenet att marknaden inte fungerar , för enbart marknadsinstrumentet leder inte till det ideala samhället .
Det är de sårbara människorna som befinner sig i det hörn där motgångarna slår .
Marknadsverkan måste användas på ett listigt sätt för att låta medborgarnas och företagens ansvar komma till sin rätt maximalt .
Om denna ansträngning misslyckas måste en statsmakt ingripa .
Kommissionens vitbok om modernisering av konkurrenspolitiken liknar mer ett diskussionsdokument .
Pläderingen för decentralisering för att lätta arbetsbördan inom Generaldirektoratet för konkurrens ger ett sympatiskt intryck , men det sätt på vilket kommissionen vill utforma denna tanke leder till att den rättsliga makten blir överbelastad .
Det går ut över rättssäkerheten för näringslivet .
Minskar verkligen kommissionens arbetsbörda när nationella domstolar är skyldiga att rapportera till kommissionen ?
Vilken åsikt har rådet om detta , och är kommissionären beredd till en grundlig omprövning av dessa punkter ?
Herr talman !
En vitbok är definitionsmässigt inte något som man tar till sig eller lämnar därhän ; den syftar till att väcka reaktioner , och det har denna vitbok helt klart lyckats med .
Den utgör ett gott diskussionsunderlag , och i den bemärkelsen är den välkommen .
Jag förstår författarnas utgångspunkter och stöder dem .
Jag utgår också från att ni , herr kommissionär , vill värna om era företrädares rykte och det de byggt upp , och att era tjänstemän har samma mål .
Jag kan inte föreställa mig att kommissionen skulle ta initiativ till att inleda en grundlig aveuropeisering eller till att börja åternationalisera .
Men jag känner ändå en viss oro , ändå har jag frågor .
För det första gäller det sammanhållningen då politiken skall omsättas i praktiken .
Allmänt sett är jag en stark förespråkare för kulturell mångfald , men inte på området konkurrenskultur på den inre marknaden .
Den inre marknaden behöver en enhetlig konkurrenspolitik , inte bara vad konceptet beträffar , utan även i fråga om att omsätta den i praktiken .
Det kommer visserligen europeiska förordningar och tolkningsmeddelanden .
Kommissionen borde också ha rätt att ta upp ärenden och ge riktlinjer åt de nationella konkurrensmyndigheterna .
Men jag ställer mig ändå frågan om vi inte löper risken att hamna i en långdragen process , där vi hela tiden skulle bli tvungna att ta ett steg tillbaka innan vi kan ta två steg framåt .
Jag skulle således vilja veta mer , herr kommissionär , om på vilket sätt kommissionen kommer att garantera en enhetlig omsättning i praktiken och om ni själv anser att de vägar som skisseras från och med punkt hundra i vitboken är genomförbara .
För det andra förstår jag näringslivets oro i fråga om rättssäkerheten .
Nu anmäls många ärenden just med tanke på detta .
I framtiden bortfaller detta instrument .
I vitboken säger ni att kommissionen ändå kommer att fatta individuella beslut som kan tjäna som riktlinjer , men vilka kriterier kommer ni att tillämpa för att den ena gången fatta ett sådant beslut och den andra gången inte ?
För det tredje vill jag gärna veta om kommissionen har undersökt vilka konsekvenser dess nya tillvägagångssätt kommer att få för näringslivets strategi .
Jag är särskilt oroad över de små och medelstora företagens öde , vilka förlorar ett visst juridiskt och ekonomiskt skydd i likhet med vad som måste vara fallet i fråga om det nya gruppundantaget för distributionssektorn .
För det fjärde skulle jag gärna vilja veta varför kommissionen inte beslutat sig för att låta nullitetssanktionen träda i kraft ex tunc då det rör sig om tydliga överträdelser av konkurrensreglerna .
För det femte handlar det om den utvidgning som står för dörren , och jag frågar mig om kandidatländerna kommer att kunna mäkta med att spela vårt spel .
I själva verket ligger de fortfarande i träning .
Vilka garantier har vi för att de kommer att växa ut till förstaklasspelare i den interna marknadens liga ?
För det sjätte och sista påminner jag om en punkt som jag också tog upp i mitt betänkande om de vertikala restriktionerna , i synnerhet företagsjuristernas så kallade legal privilege .
Om kommissionen genomför sina föresatser i vitboken förefaller det mig som om diskrimineringen på den inre marknaden mellan de externa och de interna juridiska rådgivarna kommer att bli större och således också mer oacceptabla .
Överväger kommissionen att göra något för att bevilja företagsinterna jurister i alla medlemsstater ett legal privilege ?
Herr kommissionär !
Jag ställer dessa frågor som försvarare av den inre marknaden , och jag hoppas att vi här i den bemärkelsen allesammans är partner och att diskussionen mellan dessa partner inte kommer att bli steril utan kommer att kunna bära frukt .
Herr talman !
Jag vill inleda mitt anförande om vitboken med att framföra mina gratulationer till föredragande von Wogau .
Ett tydligt bevis på den höga grad av enighet som råder mellan Europeiska socialdemokratiska partiets grupp och hans betänkande är att endast ett ändringsförslag har lagts fram under ärendets gång .
Vi ställer oss således positiva till betänkandet , precis som vi ställer oss positiva till de grundläggande inslagen i vitboken , herr kommissionär .
Gemenskapens konkurrensbestämmelser har , ända sedan fördraget trädde i kraft , varit en av gemenskapspolitikens grundvalar .
Efter nästan fyrtio år i kraft har dessa bestämmelser börjat visa sig vara föråldrade .
Därför är det angeläget med en modernisering .
Denna modernisering är nödvändig i synnerhet på fem punkter .
Punkt ett : systemet för godkännande ; punkt två : den decentraliserade tillämpningen ; punkt tre : bestämmelserna för förfarandena ; punkt fyra : rättstillämpningen och slutligen punkt fem : paragrafrytteriet .
Det har funnits ett överhängande behov av en reform av systemet för enstaka beviljanden , och en sådan har enhälligt efterfrågats av företag , forskare och advokater med specialistkompetens .
Jag har inte deltagit i en enda sammankomst för experter på gemenskapens konkurrensbestämmelser , där man inte har begärt en ändring av systemet .
Ett system som medger så pass få beslut , i form av beviljanden eller förbud , som det nu rådande systemet är inte godtagbart .
Artiklarna 81.1 och 82 har sedan länge kunnat tillämpas av de nationella konkurrensmyndigheterna .
Däremot har man inte kunnat tillämpa artikel 81.3 , något som i viss mån har förhindrat en följdriktig tillämpning av artikel 81.1 .
För närvarande har , som mina damer och herrar vet , två tyska domstolar vardera anhängiggjort ett mål för förhandsavgörande vid EG-domstolen , med ifrågasättanden av om det är möjligt att tillämpa artikel 81.1 då artikel 81.3 inte kan tillämpas .
Därför är en reform på den punkten oumbärlig .
Grunderna för konkurrensförfarandet fastslås i förordning nr 1762 .
Man röstade enhälligt för en ändring .
Det faktum att förordningen inte fastslår ett regelrätt förfarande , inte fastställer några tidsramar , inte reglerar de inblandade parternas tillgång till handlingarna och inte på ett relevant sätt erkänner rätten till försvar , har varit motiv till det enhälliga kravet på en reform .
EG-domstolen har för länge sedan godtagit att gemenskapens konkurrensbestämmelser tillämpas av medlemsstaternas rättsskipande organ , och kommissionen offentliggjorde redan 1994 ett meddelande i den frågan .
Således är det nödvändigt att underlätta ett sådant förfarande .
Paragrafrytteriet är något av det som starkast kritiseras i gemenskapens konkurrensbestämmelser .
Bedömningen av om vissa avtal är konkurrensbegränsande eller ej beror , till följd av den kontinentala rättstraditionen , snarare på en analys av avtalets klausuler än av effekten på marknaden .
Av den anledningen har det varit nödvändigt att inbegripa en ekonomisk analys .
Genom vitboken försöker man lösa dessa problem , och därför stöder vi förslagen i denna .
Vi har även upptäckt vissa brister i betänkandet .
Bland dessa kan i första hand nämnas att man , trots att det handlar om en modernisering av artiklarna 81 och 82 , lägger hela tyngdpunkten på artikel 81 och inte på artikel 82 .
I en tid då processer med samordning av företag , eller privatiseringen av monopol intar en framskjuten och till med förstärkt ställning , är det särskilt viktigt att motarbeta orimliga förfaranden .
För det andra bör förordning nr 1762 upphävas och ersättas med en ny förordning .
På den punkten stöder vi betänkandet .
Skulle däremot några av ändringsförslagen godkännas , och då i synnerhet de som framlagts av Europeiska folkpartiets grupp , anser vi att betänkandet förvanskas , att det förvandlas till ett motsägelsefullt dokument utan stringens , och i sådant fall kommer vi att bli tvungna att ompröva vårt stöd .
Herr talman , mina damer och herrar !
Bland alla de frågor som diskuteras i denna gemensamma debatt , vill jag koncentrera mig på några tankar kring det vår kollega Berenguer talade om , det vill säga den modernisering av konkurrenspolitiken som åsyftas i kommissionens vitbok .
Jag anser uppriktigt sagt att denna modernisering är tillfredsställande .
Kommissionär Monti har uppnått goda resultat i sitt arbete , precis som sin föregångare , och har tydligt visat att han , vid sidan av skapandet och utvecklandet av en inre europeisk marknad , haft förmåga att vidta de rätta åtgärderna för att marknadsekonomin inom unionen skall fungera , utan de avvikelser som vi ekonomer vet kan förekomma i samband med att marknaden expanderar , på det sätt som den har gjort inom Europeiska unionen sedan 1993 .
Om allting fungerar , om vi är nöjda , om kommissionens agerande i huvudsak har varit korrekt , varför behövs det då en ändring ?
Olika argument har lagts fram som talar för detta .
Berenguer har gjort en högst korrekt analys , där han visar på behoven och reformerna till följd av dessa i syfte att förbättra konkurrenskraften , men jag finner det angeläget att man garanterar att den standard och de kriterier som tillämpas av respektive myndighet i medlemsstaterna överensstämmer i alla avseenden .
För om de inte gör det , hamnar vi i en paradoxal situation , där kommissionen själv är den som inför illojala konkurrensmedel på den inre europeiska marknaden .
I sådana fall har vi inte gjort några framsteg , utan det skulle tvärtom innebära att vi gick bakåt i vår tillämpning av konkurrenspolitiken inom unionen .
Herr talman !
Till att börja med vill jag uttala mitt erkännande till kommissionen för den förbättring som den XXVII : e rapporten om konkurrenspolitiken i unionen innebär i förhållande till tidigare utgåvor .
Likaså vill jag framhålla det arbete som har utförts av föredragande Rapkay , som har gjort en kort och koncis analys av en så pass tjock och omfattande text som denna .
Jag stöder helt hans påpekande om behovet av att ge handlingsutrymme åt regioner - som till exempel Baskien som jag själv företräder - till följd av subsidiaritetsprincipen .
Ändå kan jag inte glömma den kritik som vid flera tillfällen har framförts , såväl av medlemsstaterna som av marknadsaktörerna som , utifrån det begränsade handlingsutrymme , den begränsade valfriheten som kommissionen har när den skall bedöma varje enskilt fall , hävdar att det rättsliga läget är osäkert , eftersom det inte finns några tydliga spelregler som gör att de inblandade kan förutse myndighetens ställningstagande och utifrån det göra korrekta ansökningar om bidrag till främjande åtgärder för den ekonomiska verksamheten och sysselsättningen , förslag om sammanslagning av bolag , etc .
Det enda säkra sättet har blivit att begära ett godkännande i förväg , via enskilda ärenden där det dröjer minst sex till åtta månader innan besked lämnas , en alldeles för lång tidsperiod som endast åtföljer problemen med bristande rörlighet till sådan verksamhet som genererar välstånd och sysselsättning .
Jag tycker att det saknas , och föreslår av den anledningen , att man fastställer ett flertal bestämmelser , tillkännager tydliga spelregler som vi alla har att vinna på : företagare , investerare , arbetstagare och befolkningen i allmänhet .
Herr talman , parlamentskolleger !
Jag vill gärna understryka att i en period av stora tekniska förändringar - se bara på det som sker inom informationstekniken eller inom andra sektorer som energi och transporter - är skyddet av konkurrensen av grundläggande betydelse för vår framtid .
När det gäller den ekonomiska tillväxten , och därmed ökningen av sysselsättning och välfärd , blir skyddet av en konkurrensfrämjande politik i våra länder inom unionen en avgörande faktor av grundläggande betydelse för vår framtid .
Det är av den anledningen jag uttrycker mitt starka stöd för den här aktuella betänkandet .
Jag har noterat att kommissionen under den senaste perioden har ansträngt sig för att hävda den principen kraftfullt och entydigt , just för att skydda marknadernas flexibilitet , såväl marknaderna för produkter som för tjänster .
Jag hävdar bestämt att detta kommer att vara av yttersta vikt för vår framtid , för den europeiska ekonomin och framför allt för att skydda vårt välstånd och den allmänna tekniska utvecklingen i Europa .
Herr talman !
För de konservativa i Storbritannien är tillämpningen av den europeiska konkurrenspolitiken på ett effektivt och enhetligt sätt kärnfrågan när det gäller att skapa en effektiv inre marknad i hela Europeiska unionen .
Därav följer att alla förslag som innebär större förändringar av systemet för att genomdriva konkurrenspolitiken måste granskas ingående och noggrant .
Sanningen är att den inre marknaden ännu inte är fullständig .
Under mina sex månader som ledamot av detta parlament har jag blivit mycket medveten om många ledamöters beslutsamhet att driva det som beskrivs som det europeiska projektet framåt .
Dagligen hör vi talas om behovet att verka för ett vidare och djupare Europa .
Men allt detta är i realiteten bara retorik när vi tittar på de nationella , regionala och lokala hinder som fortfarande står i vägen för en sann europeisk inre marknad .
Det är i detta sammanhang jag vill se kommissionens förslag .
Jag skulle vilja göra klart att vi har det största förtroende och respekt för kommissionär Monti .
Vi ser honom som mannen som skall utrota karteller .
Men han skulle förstå att vi , liksom med alla andra , måste bedöma hans enskilda förslag och underkasta dem en grundlig granskning .
Detta är vad vår föredragande i utskottet för rättsliga frågor och den inre marknaden , von Wogau , har gjort .
Jag vill gratulera honom , tråkigt nog i hans frånvaro , till det grundliga och noggranna sätt på vilket han har sammanställt detta betänkande - och också för att han har stått ut med att jag har varit så besvärlig !
Han nämnde tidigare att betänkandet antogs med en betydande majoritet , men inte med mitt stöd .
Så även om jag inte delar hans slutsatser anser jag att han i sitt betänkande har belyst många av de frågor kommissionen måste ta upp .
Den första är möjligheten att åter göra konkurrenspolitiken till en nationell fråga .
Jag vet att kommissionen är negativ till detta , men möjligheten finns .
Jag är fortfarande orolig över nationella domstolars och konkurrensmyndigheters kapacitet .
Jag är fortfarande orolig över hur den rättsliga processen som helhet fungerar .
Härom dagen frågade jag kommissionär Monti vad som händer om han har fel och konkurrenspolitiken i praktiken åter blir nationell .
Von Wogau sa att vi kan titta på EG-domstolen .
Vi i Storbritannien tittar just på EG-domstolen för tillfället .
Vi finner då att EG-domstolen inte klarar av att ge oss interimsåtgärder för en viss tvist vi har med Frankrike för ögonblicket , och där vi har kommissionens stöd .
För att ingen skall tro att detta bara är en nationell fråga tog det tio år för EG-domstolen att döma i Factortame-fallet , där den brittiska regeringen var den svarande .
Så någonting måste göras åt rättsskipningen .
Jag frågar kommissionen vad som kan göras för att snabba upp tillämpningen på detta speciella område .
Vad gäller visshet om rättsläget instämmer jag i Thyssens poäng .
Det är viktigt att företagen har visshet om rättsläget .
Jag nämnde detta för kommissionär Monti igen nyligen .
Han sade att vi inte alltid får låta oss ledas av advokater .
Jag måste säga att jag berörs av detta som advokat men också som tidigare konkurrensminister i Storbritannien .
Vi har ju alla vårt förflutna att dras med , men det är viktigt att företagen har visshet om rättsläget .
Jag skulle också vilja fråga kommissionen om den har analyserat hur denna förändring påverkar industrin : en samhällsekonomisk kostnads-intäktsanalys av det slag som nu håller på att bli en del av den europeiska politiken .
Jag vet att det har gjorts en analys av hur kommissionen påverkas av förändringen .
Vi har fått veta att människors tid slösas bort för närvarande och att förändringarna därför skulle kunna vara till fördel .
Men jag anser verkligen att vi under dessa omständigheter behöver veta vilken inverkan de får på företagen .
Slutligen söker vi som brittiska konservativa en ändrad inriktning , mot skapandet av en oberoende konkurrensmyndighet .
Jag skulle vilja höra vad kommissionär Monti har att säga om det .
Herr talman !
Alltsedan den europeiska integrationen började har Europeiska unionens konkurrenspolitik varit av central betydelse .
Den kan indelas i spänningsförhållandet , som också innefattar konceptet för den europeiska integrationen , solidariteten mellan medlemsstaterna , samarbetet mellan medlemsstaterna för att utforma bättre och mer effektiva ramvillkor för människorna och näringslivet , och konkurrensen som skall skapa impulser för att förbättra Europeiska unionens konkurrenskraft och förmåga inför framtiden .
Konkurrenspolitiken är därför med all rätt ett av de viktigaste politiska områdena .
Vi kan vara stolta över att ha en europeisk konkurrenskultur som också faktiskt syftar till att genomföra en marknadsekonomi med socialt ansvar .
Vi kan vara stolta över kartell- och fusionskontrollen .
Men vi måste vara vaksamma när det gäller de aktörer som verkar över hela världen , som det nationella agerandet inte längre kan sätta några gränser för .
Man måste tänka på en ordvändning hos den franska författaren Vivienne Forestier , som beskriver tillståndet i världen som en ekonomins terror .
Samhället överlämnar sig åt marknaden .
Så vill vi inte ha det i Europeiska unionen .
I en tidsålder av strategier rörande allianser och millenniefusioner - 1998 utbetalades 2 400 miljarder USD för övertaganden - vet vi att en konkurrensskadlig praxis stävjas inte bara med hjälp av våra egna bestämmelser , utan också via bilateralt samarbete med USA eller Japan eller andra , så länge det fortfarande inte finns någon internationell konkurrensrätt , som absolut borde finnas !
Europeisk konkurrenspolitik - detta glömmer vi ofta bort - är inte bara av betydelse för den rättvisa konkurrensen som sådan , utan också för prisutvecklingen , tillväxten och sysselsättningen och därmed också för medborgarna .
Liksom de andra kollegerna kräver jag medbeslutande från Europaparlamentet när det gäller konkurrensrätten .
Det måste äntligen genomföras !
Det är också viktigt att framhäva sammanhanget mellan konkurrenspolitik och konsumentskydd .
Det är positivt att kommissionär Monti på detta område vill uppnå framsteg i dialogen med Europaparlamentet , men också i dialogen med de icke-statliga organisationerna , konsumentskyddsorganisationerna och medborgarna .
Större öppenhet kommer också att bidra till en offentlig acceptans av konkurrenspolitiska beslut .
Då kan man nämligen förstå , att exempelvis de lägre el- och telekommunikationspriserna också är ett resultat av den europeiska konkurrenspolitiken och att Bryssel inte bara måste ställas vid skampålen när det fattas beslut om stöd , som i en aktuell eller lokal situation säkert kan förorsaka problem .
Det måste också finnas klarhet särskilt om konkurrensreglerna med tanke på utvidgningen av EU .
Det måste då framhävas att en statlig stödpolitik - detta framgår också tydligt av Jonckheers betänkande - även i fortsättningen måste ge varje stat friheten att självständigt definiera och utforma sina offentliga uppgifter och ägandeförhållanden .
Det måste därvid stå klart att stöden kan ha en nyttig funktion för att utjämna misslyckanden på marknaden och främja gemenskapens mål .
Ett påpekande om vitboken : Revideringen av artiklarna 81 och 82 innebär en vändpunkt i fråga om kartellbestämmelserna .
Jag vänder mig mot detta , i motsats till majoriteten i denna kammare och även till majoriteten i min egen grupp , eftersom jag anser att systemet med direkt tillämplighet av undantagsregeln konkurrenspolitiskt är klart underlägset ett system där man har förbud med administrativt förbehåll , och därför att jag ser risken för en åternationalisering .
Det rådande systemet medger öppenhet och erbjuder rättssäkerhet för företagen ; dess anmälningsplikt har utan tvivel lett till disciplinering och avskräckning .
Problemet med för stor arbetsbörda som av kommissionen ställs i förgrunden är inte någon tillräcklig anledning till en djupgående ändring av rättssystemet .
Här måste man också fråga sig om det över huvud taget kan genomföras utan en ändring i fördraget .
Herr talman !
Jag är mycket glad att Randzio-Plath nämnde den mycket viktiga bakgrunden till vår debatt , eftersom ingen talare hittills har gjort det .
Eurons tillkomst i början av förra året släppte lös en enorm konkurrenskraft inom den europeiska industrin vilken bemöts av en sammanslagningsvåg av aldrig tidigare skådade proportioner .
Till exempel visar nu siffrorna för förra året att det totala värdet av fusioner inom Europa var 1,4 triljoner euro , vilket är sju gånger så mycket som vid höjdpunkten för den senaste europeiska fusionshaussen 1990 .
Detta ställer konkurrenspolitiken inför enorma utmaningar , vilka jag hoppas att den kommer att leva upp till , eftersom många av dessa sammanslagningar helt visst kommer att vara utformade för att skydda företagens vinstmarginaler mot konkurrens snarare än att enbart stärka produktiviteten och ge dessa företag förmåga att verka i större skala .
Kommissionär Monti och hans kolleger står inför en ofantlig utmaning och ELDR-gruppen är angelägen om att konkurrenspolitikens framstötar inte försvagas vare sig vad gäller granskningen av fusioner eller övervakningen av kartell- och monopolfrågor .
Visst kan man delegera till nationella myndigheter , men vi skulle då vilja betona vad von Wogau sade i sitt betänkande om behovet av en regelbunden övervakning av de nationella myndigheterna för att se till att det europeiska maskineriet inte slirar och speciellt be kommissionären att försäkra oss om att det dessutom kommer att förekomma stickprovskontroller .
Herr talman !
Jag vill under den korta talartid som står till mitt förfogande uttala mitt stöd för det arbete som har lagts ned av samtliga föredragande och även stödja mycket av det som här har sagts , i synnerhet av min kollega Jonckheer , som kritiserar den alltför omfattande sammanställningen av fakta och påpekar behovet av insyn och av en socioekonomisk balans vad stödet beträffar .
Jag delar även kritiken mot att inget avseende har fästs vid artikel 82 , framför allt med tanke på att vi kan tillgripa oriktiga metoder vid en koncentration av marknaden .
I egenskap av ledamot från Baskien , vill jag uttala mitt fulla stöd för åtgärder som att tillämpa en vederbörlig konkurrens på marknaden .
Jag vill påpeka detta om det nu skulle råda några tvivel angående den kritik vi riktat mot kommissionen i allmänhet och mot Monti i synnerhet , på grund av dennes attack mot stimulansåtgärderna till de baskiska företagen och det faktum att han betraktar dessa som ett statligt stöd .
Det vi skulle reagera negativt på är om kommissionen gick vidare utan att ha förstått det inre väsendet hos det generella systemet i vår ordning , med ett medansvar , som innebär att våra baskiska taxeringsnormer är av samma karaktär , att grundsatserna och målsättningen med dessa är samma som för normerna i unionens stater , och att dessa normer gäller alla skattebetalare som på ett eller annat vis omfattas av dem .
Herr talman , herr kommissionär !
Ja , vi behöver konkurrens !
Vi behöver konkurrens för att få så låg arbetslöshet som möjlighet , för att få en välutvecklad hälsovård , social rättvisa , hög social standard , och vi behöver naturligtvis också - det är nationalekonomiska konkurrenskriterier - en företagsekonomisk konkurrens : högsta kvalitet på produkterna , samma villkor för tillgången till marknaden för alla företag , miljövänliga produkter .
Det betyder att vi måste lyckas koppla samman de nationalekonomiskt erforderliga konkurrenskriterierna med de företagsekonomiska .
Jag får ofta intrycket att i motsats till hur det förhöll sig i det land som jag kommer från - Östtyskland - där den nationalekonomiska konkurrenskraften var närmast allenarådande och den företagsekonomiska inte beaktades , gör man nu ofta motsatsen ; samhället tänker nästan enbart företagsekonomiskt .
Detta säger jag själv som företagare , som absolut är intresserad av detta .
Men på det viset kan ett system inte fungera !
Det måste finnas en koppling .
Jag vill ge er ett exempel : Europeiska unionen har med all rätt stött stålverket Grönitz i Brandenburg , fastän endast 700 arbetstillfällen återstår av 5 000 .
Men det är konkurrenskraftiga arbetstillfällen , ty detta stålverk är nu nummer 2 bland verktygsstålstillverkarna i Förbundsrepubliken Tyskland .
Den som nu i princip äventyrar produktionen i detta stålverk genom att kräva tillbaka det tidigare godkända stödet , äventyrar inte bara själva stålverket , utan han äventyrar i denna region en arbetsgivare som naturligtvis även små och medelstora företag är beroende av .
Detta kan naturligtvis inte vara Europeiska unionens konkurrenspolitik !
Om vi vill ha konkurrens , då måste vi få till stånd denna koppling mellan de nationalekonomiska nödvändigheterna och de företagsekonomiska förutsättningarna .
Det är också den enda chansen att bygga upp regionala ekonomiska kretslopp i de underutvecklade regionerna på detta sätt , som innebär att det finns en social trygghet för människorna och att köpkraften stärks .
Därmed måste vi också ta avsevärt mycket större hänsyn till en ekonomisk politik som är inriktad på efterfrågan , än till en som är enbart utbudsinriktad .
Herr talman !
Inte sedan jag valdes in i detta parlament 1994 har jag sett ett betänkande med så anti-irländska känslor och övertoner som Jonckheers betänkande som vi diskuterar i dag .
Jag skulle vilja citera betänkandet ord för ord : " Det statliga stödet per capita är störst i Italien , Tyskland och Irland .
Irland är dock det land som får mest stöd om man lägger ihop det nationella stödet och gemenskapens regionala och sociala stöd . "
Jag anser att föredraganden bara leker med siffror .
Jag har svårt att inse hur han kan stoppa in regionala och sociala fonder i denna matematiska ekvation .
Jag skulle vilja påminna ledamoten om att Europeiska unionen har antagit de nya riktlinjerna för regionalstöd för perioden efter år 2000 .
Detta var bara en förlängning av de politiska målsättningarna att komplettera den inre marknaden i Europa .
Regionala skillnader måste övervinnas om den inre marknaden skall lyckas och frodas .
Det faktum att ett stöd på 40 procent med ytterligare 15 procent till små och medelstora företags fasta investeringskostnader kommer att beviljas för företag som startas i mål 1-regioner i Europa efter år 2000 är välkommet .
Jag påminner Jonckheer om att irländska företag och utländska företag i Irland fortfarande måste ta sig över två hav för att komma till marknaden på det europeiska fastlandet .
Ingen annan medlemsstat har ett så ogynnsamt läge .
Herr talman , mina damer och herrar , kära kolleger !
Kartellförbudet utgör kärnan i en fungerande konkurrensordning i Europa .
Det praktiska hanteringen av övervakningen av kartellförbudet har kommissionen funnit vara otillfredsställande ; det kan man till att börja med hålla med om .
Men i fråga om lösningen skiljer sig åsikterna åt .
Kommissionens förslag avviker formellt inte från kartellförbudet , men till sitt resultat är detta förslag en övergång från ett förbud med godkännandeförbehåll till ett godkännande med förbudsförbehåll .
Detta är en växling från förbudsprincipen till missbruksprincipen .
En så graverande systemändring avvisas beslutsamt av mig och andra kolleger .
Jag godtar inte att ett problem med det praktiska genomförandet skall ge anledning till att ändra rättsordningen .
Vi ändrar på rätten för att det åter skall gå att verkställa den ; det anser jag inte vara godtagbart .
Kommissionen avstår från sitt monopol att ge undantag för vissa slag av stöd .
Mot bakgrund av detta planerade system med direkt tillämplighet av undantagsregeln är konkurrensbegränsningar utan vidare undantagna , såvida det föreligger förutsättningar enligt artikel 81.3 EG-fördraget .
Nödvändigheten av anmälningar till Bryssel faller bort , vilket innebär att kommissionen i denna sak kommer att flyga med autopilot i framtiden .
Det finner jag inte godtagbart .
Kommissionens koncept kompletteras genom en ökad kontroll i efterhand av de nationella myndigheterna och domstolarna i medlemsstaterna .
Här kommer vi emellertid , om det äger rum på detta vis inom ramen för en åternationalisering , att få en konkurrenspolitisk trasmatta i Europa .
Jag tror inte det är godtagbart .
Här försvagas en kärnpunkt i den europeiska politiken .
Den av kommissionen planerade systemändringen i den europeiska kartellrätten är konkurrenspolitiskt sett synnerligen riskabel .
Vi har tillräckligt med andra optioner i det befintliga systemet för att säkra öppna marknader och fri konkurrens .
För övrigt kommer kommissionen med sitt förslag åter tillbaka till gamla förslag , som lades fram redan någon gång på 50- och 60-talet .
De fick ingen majoritet .
Eftersom Frankrike då mycket starkt ställde undantagsregeln i förgrunden , kompenserades man av eftergifter inom jordbrukspolitiken .
Fyrtio år senare dyker detta förslag nu upp igen , och det kommer - det är jag säker på - att ge utrymme för kartellbildningar till nackdel för konsumenterna i Europa .
Jag anser inte att det är godtagbart !
Herr talman , kära kolleger !
I denna viktiga konkurrensdebatt vill jag i dag mera särskilt uttala mig om Langens text , om gemenskapens regler för stöd till stålindustrin .
Stålsektorn är särskilt känslig för konkurrensstörningar , något som EG-domstolen erkände år 1996 .
Jag drog för övrigt själv samma slutsats för några år sedan , i ett betänkande om den europeiska stålindustrins styrka och svaghet .
Det var därför berättigat att inrätta ett stödsystem för denna sektor , i syfte att garantera de livskraftiga företagens överlevnad , även om det stod i strid med artikel 4 i EKSG-fördraget .
Detta är syftet med den sjätte regeln för stöd till stålindustrin .
Men samtidigt är det viktigt att förhindra att konkurrensvillkoren kränks och att marknaden utsätts för allvarliga störningar , därav vikten av att fastställa regler för den här typen av stöd .
Det är således nödvändigt att även i fortsättningen begränsa statsstöden till följande områden : forskning , utveckling , miljöskydd samt nedläggningar av företag .
Av samma skäl är det ytterst viktigt att medlemsstaterna uppfyller förpliktelsen att till kommissionen anmäla de stöd som de beviljar sina stålföretag .
Kommissionen föreslår snävare tidsramar .
Jag instämmer i det förslaget .
I likhet med föredraganden gläder jag mig åt kommissionens rapport , men beklagar ändå att den inte täcker alla aspekter av dessa stöd .
Trots att gemenskapens regler om stöd till stålindustrin formuleras på ett mycket tydligt sätt , har kommissionen beviljat stöd till stålföretag som inte tillhör någon av de kategorier som åsyftas i reglerna .
Med omsorg om rättvisa bör man antingen tillämpa reglerna eller ändra på dem .
För att till sist avsluta , herr talman , krävs det en översyn av reglerna innan EKSG-fördraget löper ut , för jag anser att stödsystemet bör finnas kvar efter år 2002 .
Jag är följaktligen positiv till att en förordning från rådet skall erbjuda en garanti i det avseendet .
Därför väntar vi - jag inväntar förslag från Europeiska kommissionen med den innebörden .
Herr talman !
Även jag kommer att tala om Langens betänkande beträffande stödet till stålindustrin .
Jag håller med föredraganden på två punkter .
För det första vad gäller behovet av att garantera lika villkor för stödet till alla medlemsstater , och för det andra vad gäller stödets genomblickbarhet .
Vi kritiserar , precis som föredraganden , att kommissionen trots de normer som härrör sig från det sjätte regelverket om stöd till stålindustrin , vid flera tillfällen har beviljat stöd till företag som inte överensstämmer med kategorierna för reglerna .
Hur som helst , herr talman , det som mest bekymrar oss är sänkningen av priserna med 30 procent till följd av importen .
Orsaken till denna prissänkning är den illojala konkurrensen från Sydkorea och Taiwan inom stålindustrin , på grund av andra villkor för arbete och stöd .
Orderingången inom stålindustrin och sjöfartssektorn - den frågan diskuterade vi nyligen - har minskat drastiskt med en minskad sysselsättning som följd .
Jag bor i en region där sjöfartssektorn för närvarande lider av stora problem : Asturien .
För marknader med internationell räckvidd bör det finnas arbetsnormer med internationell räckvidd och stöd med internationell räckvidd .
Jag vet att det är svårt att åstadkomma något sådant nu , men om vi inte lyckas åstadkomma rättvisa arbetsnormer för alla arbetstagare , både här och i övriga världen , om vi inte kan åstadkomma ett rättvist stöd för alla länder , både här och i övriga världen , kommer det att bli mycket svårt att bibehålla sysselsättningen , både i Europa och i övriga världen .
Herr talman , herr kommissionär , herr generaldirektör , mina damer och herrar !
Jag vill framför allt konstatera följande beträffande von Wogaus betänkande : Jag välkomnar kommissionens ansträngningar att utan något tabu inleda en diskussionsprocess om de hittills benhårda reglerna om förfarandena , och föreslå konkreta reformåtgärder .
Jag gratulerar föredraganden Karl von Wogau , som tar itu med saken , men också helt konkret kräver klargöranden , hänvisar till erforderliga åtföljande åtgärder och kritiskt kallar de aktuella uttalade problemen vid deras rätta namn .
Vitboken och betänkandet bidrar i inledningsskedet till en process av nödvändig eftertanke , nödvändiga diskussioner och reformer , som ännu inte är avslutad , eftersom somliga frågor fortfarande måste redas ut av oss , av domarna , medlemsstaterna och framför allt av de berörda små och medelstora företagen .
Konkurrenspolitiken måste även i fortsättningen hanteras centralt och kommer inte att åternationaliseras , eftersom detta skulle äventyra den inre marknaden och handelsplatsen Europa i den globala världsekonomin .
Men den måste europeiseras på ett sätt som motsvarar subsidiariteten .
Jag välkomnar därför också att ansvaret läggs på den enskilde , utan att kommissionen undandrar sig sitt ansvar .
Erfarenheterna i praktiken - endast 9 fall avvisades , och 94 procent av de fall som kommissionen skulle bearbeta klarades av inte formellt , utan endast med hjälp av icke offentliggjorda , rättsligt icke bindande administrativa skrivelser eller helt enkelt på grund av att tiden gick - visar tydligt att man måste sätta tidsmässiga , personella och finansiella gränser för kommissionens arbete i en tidsålder av globalisering och EU-utvidgning .
Avslutningsvis vill jag säga vad jag förväntar mig av denna reform : en rättvis konkurrens och lika konkurrensvillkor , rättssäkerhet för alla företag , en enhetlig tillämpning av konkurrenspolitiken , förenklade förfaranden enligt principen one-stop-shop , en samordning av de nationella och för mig oberoende konkurrensmyndigheterna , ett nära samarbete mellan de nationella myndigheterna och domstolarna och kommissionen , liksom en klar ansvarsfördelning mellan nationella myndigheter och domstolar vid tillämpningen av den europeiska konkurrens- och kartellrätten ; av kommissionen förväntar jag mig att den koncentrerar sig på väsentligheterna genom att fullgöra sina uppgifter som högsta väktare av den europeiska konkurrenspolitiken .
Jag väntar med spänning på att få se hur diskussionerna , som förs på bred basis , kommer att mynna ut i det första lagförslaget .
Kommissionens rapport bekräftar att de statliga företagsstöden ökar , Tyskland undantaget .
Men det enda som oroar kommissionen är konkurrensvillkoren .
Vi sätter oss däremot in i arbetarklassens intressen .
Samhället tjänar ingenting på de enorma överföringarna av offentliga medel till privata företag .
Titta på bilbranschen ; där har statliga subventioner och olika former av statsstöd ökat med 24 procent under den granskade perioden .
Av vilka skäl då ?
Inte för att bevara arbetstillfällen .
Alla dessa företag har avvecklat arbetstillfällen , ja t.o.m. avskedat folk .
Och det är inte för att förbättra arbetsvillkoren , för arbetsvillkoren försämras när färre arbetare skall producera mer .
Var dessa företag i behov av statliga stöd för att överleva ?
Nej , biltillverkarna håvar in kolossala vinster sedan flera år tillbaka .
De statliga stöden får inte endast negativa bieffekter då de främjar en jakt på subventioner genom omlokaliseringar från ett land till ett annat , vilket medges i Jonckheerbetänkandet ; de är också oacceptabla eftersom de innebär att offentliga medel används för att berika en handfull privata aktieägare .
Eftersom man överallt gynnar de rikaste med hjälp av statens pengar , inskränker man också det sociala skyddet överallt i Europa - man överger den offentliga sektorn , man lägger ner sjukhus .
Genom att rösta emot Jonckheerbetänkandet vill jag hävda att det krävs en annan politik , dvs. att alla stöd till privata företag stoppas och att de därmed frigjorda pengarna används för att utveckla tjänster av allmänt intresse och för att anställa personal inom den offentliga sektorn .
Herr talman !
Dagens debatt är utomordentligt viktig , för konkurrensprincipen har förmodligen varit hörnstenen för den inre marknaden .
Som ett sätt att tillämpa konkurrensprincipen har man utformat artiklarna 85 till 94 , konkurrenspolitiken närmare bestämt , granskningar av sådant statligt stöd och sådana skattebestämmelser som skulle kunna förändra konkurrensen .
Till en början de indirekta skattebestämmelserna ; och nyligen , tack vare kommissionär Monti , de direkta bestämmelserna , och då i synnerhet uppförandekoden .
Detta har fungerat tämligen väl , men tiden går , precis som i den välkända filmen Casablanca , och det är nödvändigt att anpassa de bestämmelser som vi hittills har tillämpat till de nya omständigheterna .
Jag har lagt märke till en stark enighet på den punkten i alla anföranden .
För det första är det nödvändigt att man i utformningen av bestämmelserna gör upp tydliga och heltäckande regler .
Förmodligen är förekomsten av oklara regler , oreglerade områden eller regler som endast fastslår vaga juridiska begrepp allvarligare i denna del av bestämmelserna än i andra delar .
Inte minst - så som fallet är i reformens andra del - då tillämpningen av bestämmelserna överlåts åt de nationella myndigheterna .
För det tredje , anser jag att kommissionen har en viktig roll att fylla i och med att man motstår frestelsen att inrätta oberoende byråer , något som skulle förändra kommissionens innersta väsen , som ett sätt att garantera en enhetlig tillämpning från de internationella organens sida .
Och slutligen för det fjärde- och det har redan påtalats - har den internationella rättsordningen förändrats .
Det kunde vi se i och med den misslyckade konferensen i Seattle och nu ser vi det i samband med de bilatera konferenserna för olika regioner eller länder .
Konkurrensprincipen bör ha en universell tillämpning .
Och vi bör se till att miljönormerna , arbetsnormerna följs , för att undvika dumpning på det området , att rätten till egendom respekteras fullt ut , att det sker en granskning av det statliga stöd som - precis som det har sagts här - snedvrider konkurrensen inom flera sektorer och förstör sysselsättningen på hemmaplan , och vi bör definitivt se till att snarlika villkor tillämpas som förhindrar att stödåtgärder , snedvridningar på den inre marknaden i andra länder sprids till internationell nivå genom fusk .
Herr talman , herr kommissionär Monti !
Jonckheers betänkande om statliga stöd till tillverkningsindustrin och vissa andra sektorer innehåller mycket gott .
För det första framhåller man i betänkandet parlamentets fasta ståndpunkt att de statliga stöden målmedvetet måste minskas för att den inre marknaden skall kunna fungera korrekt .
Många av betänkandets slutsatser vållar dock åtminstone inom vår grupp allvarlig oro .
Att sådana här översikter är nödvändiga bevisas till exempel av det faktum att mängden av och nivån på det statliga stödet per capita varierar kraftigt mellan olika medlemsstater .
Stöd som väller fram till följd av nationella egoistiska utgångspunkter ger företagen orättvisa fördelar , snedvrider på det sättet konkurrensen och leder till en ineffektiv och oekonomisk fördelning av de knappa europeiska resurserna .
Det är inte heller helt oväsentligt vilka typer av stöd det handlar om .
Statliga stöd som förutsätter egna ansträngningar av stödmottagaren måste prioriteras .
De statliga garantierna till exempel , angående vilka kommissionen nyligen offentliggjort ett ställningstagande , måste naturligtvis räknas till de statliga stöden men är enligt min mening ett bättre alternativ än direkta bidrag till företag .
Rapporten om konkurrenspolitiken framhäver vidare kommissionens tro på kraftig reglering i stället för att betona de ekonomiska effektivitetsargument som påverkar konkurrenskraften .
Den europeiska ekonomin kommer aldrig att uppnå önskad konkurrenskraft om vi inte visar att vi litar på marknadens funktion .
Om konkurrenspolitiken skall underordnas social- och miljöpolitiska ambitioner kan vi bara drömma om verklig effektivitet och ekonomisk tillväxt .
Konkurrenspolitiken måste också ses som en del av den ekonomiska helheten och den måste bedömas bland annat i förhållande till handelspolitik och immateriella rättigheter .
Man kan inte enbart betona dess sociala dimension .
Socialpolitiska mål uppnås bäst genom en kraftigare ekonomisk tillväxt , inte genom att kompromissa om konkurrenspolitiska lösningar .
I Rapkays betänkande betonas också konkurrensrättens internationella dimension .
Jag tycker också att det är bra om man på internationell nivå uppnår samförstånd när det gäller vissa konkurrensrättsliga kärnprinciper .
Om man däremot strävar efter enhetliga miniminormer leder detta lätt till att man går den enklaste vägen och väljer den minsta gemensamma nämnaren , vilket urvattnar alla konkurrenspolitiska mål .
Herr talman , kommissionär Monti !
Uppdateringen av konkurrensreglerna borde vara en viktig uppgift för Europeiska unionen , inte bara mot bakgrund av och som en konsekvens av de förändringar som inträffat genom åren , utan också med tanke på unionens förestående utvidgning .
Jag tackar föredraganden Karl von Wogau för det engagemang han lagt ner och jag uppskattar verkligen hans resonemang .
Jag vill också uttrycka min uppskattning för de synpunkter som jag har fått från professor Tesauro , ordförande för den italienska myndigheten , och som jag är övertygad om att professor Monti i en anda av samförstånd kommer att ta vederbörlig hänsyn till .
Det problem vi står inför är utan tvekan hur vi skall kunna ytterligare avreglera marknaden och framför allt se till att de olika nationella marknaderna blir homogena , de marknader som för tillfället uppvisar stora skillnader , skillnader som tydligt framkommer om man jämför den engelska marknaden med den italienska och franska .
På den senare finns det starka inslag av statlig protektionism , något som inte finns på den engelska och som är ytterligt begränsat i Italien .
Ett annat problem är ekonomierna i de länder som berörs av utvidgningen , som riskerar att för evigt bli subventionerade ekonomier om det inte kan ske en gradvis anpassning .
Enligt min mening är det även nödvändigt att skapa en nivå där man skall införa två viktiga inslag som karakteriserar vårt ekonomiska system : de små och medelstora företagen , som utgör det sammanbindande elementet i den europeiska ekonomiska verkligheten , och det sociala skydd som Europa alltid har garanterat de ekonomiskt svagaste grupperna .
Skyddet av marknadens sociala dimension utgör hela skillnaden mellan en total marknadsliberalism och ett system som skall kunna förbättra människors livskvalitet .
En aspekt som måste beaktas i det nya regelverket utgörs av ekonomierna i de ultraperifera regionerna och i öregionerna , som behöver skyddas .
Därför tror jag att det skulle vara lämpligt att även tänka på att skapa två fokus för den externa marknaden och att inleda ett givande samarbete med Ryssland och Medelhavsländerna , just för att de ekonomierna skall bli mindre perifera .
Jag hoppas - och i det sammanhanget vill jag tacka professor Monti - att man i det nya regelverket ägnar ett så stort utrymme som möjligt åt den ekonomiska politiken och att man verkligen garanterar dess sociala funktion .
Herr talman !
Konkurrens är hjärtat och kraften i den europeiska politiken för den inre marknaden .
En fri öppen marknad kan bara existera under konkurrensens överhöghet , begränsad av tydliga , enhetliga spelregler .
Karl von Wogau förordar detta på ett mycket bra sätt i sitt betänkande .
Men Europa förändras .
Ekonomierna växer , vi expanderar till 25 till 30 medlemsstarter .
Europeiska kommissionen kommer att bli överbelastad om den nuvarande politiken skall fortsätta .
Det är därför nödvändigt med en modernisering av konkurrenspolitiken .
Det råder ingen diskussion om detta .
Men trots detta kan jag ändå inte släppa en oro i fråga om den planerade decentraliseringen .
På vilket sätt kommer kommissionen som fördragens väktare att garantera att man på ett enhetligt sätt fattar beslut i konkurrensärenden i London , Palermo , Helsingfors och inom kort i Budapest och Ankara ?
Det är nödvändigt att förhindra olikhet inför lagen , annars skulle en strid ström av konkurrensmål gå till den domstol där den mildaste bedömningen görs .
Det räcker inte med att säga att medlemsstaterna redan har 40 års erfarenhet .
I Nederländerna ligger konkurrensmyndigheten fortfarande i sin linda .
Detta land har att göra med en mycket liten marknad som tyvärr ofta samtidigt definieras som den relevanta marknaden .
Detta i motsats till Tyskland , där en mycket erfaren Kartellamt utövar sina befogenheter på en gigantisk marknad .
Europeiska kommissionens tilltro till att tolkningen av lagstiftningen kommer att vara lika i alla väderstreck är vad vi i katolska kretsar kallar " övermodigt förtroende " , och det är förbjudet .
Det krävs mer arbete för att uppnå enhetlighet .
Jag tänker på specialiserade , nationella domstolar med möjlighet att överklaga direkt till en särskild konkurrensdomstol vid EG-domstolen .
Denna särskilda domstol behövs på grund av att det är nödvändigt att bygga upp en bred expertis .
Dessutom tillåter inte de mycket stora ekonomiska och sociala intressen som hör samman med ärenden av den arten att ett domslut låter vänta på sig i två år , vilket nu är helt normalt .
Vad anser kommissionären om detta ?
Jag vill avsluta med en viktig punkt för det lilla och medelstora företaget .
För att skapa trygghet för det lilla och medelstora företaget bör Europeiska kommissionen själv utarbeta en undantagsförordning för det lilla och medelstora företaget i syfte att också möjliggöra horisontala undantag vid sidan av vertikala .
Småföretagare måste genom samarbete kunna försvara sig mot de stora kedjorna .
Syftet med den europeiska konkurrenspolitiken kan inte vara att göra livet omöjligt för småföretag .
Vad småföretag beträffar bör man dessutom begrunda om det inte skulle kunna vara lättare att hantera ett system med en varning i förväg , gult kort , i stället för att omedelbart ge ett rött kort som kommer att fungera som böter och hota företagets fortlevnad .
Herr talman !
I egenskap av sista talare har jag privilegiet , herr kommissionär , att få tala om att majoriteten av den här församlingen stöder ert initiativ och har visat ett fullständigt , och jag tror även högst berättigat förtroende för er som kapten på den här skutan .
Men vi vill utgöra besättningen på skutan , eftersom vi befinner oss på samma skuta som ni .
Därför anser jag att en interinstitutionell dialog är oumbärlig , så att vi kan precisera och nyansera denna så viktiga reform och föra den i hamn .
De förslag som har lagts fram här kan delas in i tre stora grupper .
I första gruppen finns den oro som vissa av oss har gett uttryck för , och då i synnerhet Randzio-Plath , ordförande i utskottet för ekonomi och valutafrågor , en oro för att detta nya system som ett rättsligt undantag inte skall överensstämma med fördraget .
Jag delar hennes oro och anser att den saken bör undersökas .
I andra gruppen ingår frågan om företagens rättssäkerhet .
Det är sant , herr kommissionär , att kommissionen inte är en maskin som tillverkar rättssäkerhet .
Det kan vi alla vara överens om .
Men det är likaså sant - och det har alla sektorer i den här församlingen upprepat - att den europeiska industriella vävnaden är en vävnad som består av små och medelstora företag , och att kommissionen många gånger är den som företräder auctoritas , legitimering , legitimitet , av det som är den inre marknaden .
På den punkten vill jag framföra min åsikt om något Karas sade .
Det har endast förekommit nio beslut om avslag .
Där har jag nytta av min erfarenhet som advokat .
Hur många gånger har det inte hänt att en advokat med två bolag och ett projekt har ändrat projektet efter en orientering ex ante från kommissionens sida , för att det skall överensstämma med konkurrensbestämmelserna !
Det är därför en aspekt att ta hänsyn till .
I den tredje gruppen ingår problemet med en enhetlig tillämpning av gemenskapsrätten .
Thyssens utmärkta inlägg kunde knappast ha varit bättre .
Jag anser att det är bra med ett biologiskt mångfald , och även med ett kulturellt mångfald , däremot inte med ett mångfaldigt tillämpande av rätten , av det som är själva kärnan i den inre marknaden , det vill säga , konkurrensbestämmelserna .
Där krävs en närmare precisering .
Endast i vissa länder , som i Tyskland , har man en specialiserad rättsskipning .
Måhända är det en lösning som är värd att undersöka , men vi bör även undersöka andra möjligheter .
Det vi inte får göra , herr kommissionär - och med detta vill jag avrunda - är att ge så mycket som ett lillfinger , och än mindre räcka vapen åt dem som talar om de europeiska institutionerna som en fråga för de mäktiga , för de inflytelserika , för de rika , och inte för den enskilda medborgaren , inte för de små och mellanstora företagen , som skulle känna sig utelämnade åt sina värsta föreställningar- som aldrig kommer att förverkligas , för de rätta åtgärderna kommer att vidtas för att undvika något sådant - till domstolar som avkunnar olika domar , mycket sent , utan några realistiska möjligheter till kontroll annat än med det som fransmännen kallar le parcours du combattant , det vill säga efter jag vet inte hur många år , när domstolen i Luxemburg uttalar sig , en domstol som vi alla vet för närvarande är starkt överbelastad .
Herr kommissionär , vi står inför en reform som jag inte nog kan poängtera vikten av .
Effekten av denna reform sprider sig till konkurrensen , den sprider sig till sammanhållningen på den inre marknaden , jag tror att den på djupet påverkar det som är meningen med den europeiska integrationen , meningen med den europeiska integrationens legitimitet .
Därför , herr kommissionär , räknar vi med denna interinstitutionella dialog som ett sätt att närmare precisera en reform som vi alla hoppas och tror att vi kommer att ro i hamn med er som kapten och oss som besättning .
Herr talman , ärade ledamöter !
Låt mig varmt tacka utskottet för ekonomi och valutafrågor och hela Europaparlamentet för det stora intresse de visar för konkurrensfrågorna .
Denna gemensamma debatt är , herr talman , enligt min åsikt ett levande och starkt bevis på detta .
Vi har lyssnat på resonemang av stor djupsinnighet som samtidigt har rört ekonomisk politisk filosofi och institutionernas arbete .
Vår gemensamma avsikt är att uppdatera , förstärka konkurrenspolitiken , grundbulten i den sociala marknadsekonomin och det europeiska konstruktionsarbetet .
Den röda tråden i arbetet med att reformera konkurrenspolitiken , som vi skall genomföra gemensamt , är syftet att garantera ett säkrare skydd för konkurrensen , minska den byråkratiska börda som tynger företagen , och att föra beslutsprocesserna närmare medborgarna .
Jag vill personligen varmt tacka von Wogau för det engagemang han visat i arbetet med vitboken och för den goda kvaliteten i hans betänkande .
Låt mig sammanfatta de synpunkter som framförts i debatten om von Wogaus betänkande i fyra punkter , som jag inte anser vara kritik mot kommissionen , utan snarare som bidrag av avgörande betydelse , eftersom det finns invändningar som det är viktigt att framföra och som vi tillsammans vill reda ut : frågan om effektiviteten , frågan om risken för åternationalisering , frågan om en enhetlig tillämpning , frågan om rättssäkerheten .
Låt mig som hastigast gå igenom dem en efter en .
Effektiviteten : jag är övertygad om att denna reform kommer att göra det möjligt för oss att förstärka , snarare än försvaga , konkurrensskyddet inom ramen för den inre marknaden .
Det nuvarande anmälningssystemet , ärade parlamentsledamöter , tillåter oss inte längre att uppnå det målet eftersom det inte garanterar information till kommissionen om de allvarligaste restriktionerna - låt mig påminna om att under trettiofem år har endast nio beslut om förbud fattas som en följd av en anmälan och där det har saknats en stämning - inte garanterar öppenhet och inte medför en reell rättssäkerhet för företagen som , i de flesta fall , mottar ett enkelt administrativt meddelande som sedan arkiveras .
Det system som föreslås gör det möjligt att förbättra konkurrensskyddet , framför allt därför att det kommer att tillåta kommissionen att koncentrera sin uppmärksamhet på de allvarligare inskränkningarna , just därför att det i högre grad kommer att engagera de nationella konkurrensverken i arbetet att hålla nere kränkningarna och , slutligen , för att det gör det möjligt för dem som drabbas av kränkningarna att vända sig direkt till de nationella rättsinstanserna , vilkas uppgift det är att skydda de enskildas rättigheter .
Frågan om åternationaliseringen : först av allt , även om det skulle vara överflödigt , skulle jag vilja påminna om och understryka , tre gånger om det är möjligt , att vitboken inte i något avseende berör frågan om koncentrationer och statliga stöd - vi överväger inte en tillbakagång i det avseendet - utan , när det gäller förordning 17 , så finns det en risk för åternationalisering .
Ni kan föreställa er att vi naturligtvis har ställt oss den här frågan : vi har ställt oss frågan och vi följer den uppmärksamt , även tack vare den oro som ni har givit uttryck för .
Men jag tror uppriktigt sagt inte att denna oro är berättigad .
Kommissionens förslag ger kommissionen en central roll när det gäller att bestämma konkurrenspolitikens inriktning .
Reformen innebär ingen minskning i kommissionens verksamhet , utan en koncentration av uppmärksamheten till de viktigaste fallen .
Reformen kommer att leda till en gradvis utveckling låt mig understryka detta för jag tyckte om den formulering som användes av ordföranden Randzio-Plath och som jag för övrigt helt instämmer i - av en europeisk konkurrenspolitik .
Reformen kommer att leda till en överföring , en omplantering på den europeiska konkurrenskulturens mark - där det i dag växer diverse olika plantor , som verkligen inte är enhetliga - av de olika nationella konkurrenskulturerna .
Det kommer att leda till att man gradvis överger de femton olika nationella rättssystemen till förmån för en vidare tillämpning av gemenskapsrätten , som kommer att kunna tillämpas av allt fler aktörer .
Detta , tillåt mig understryka det , är att göra konkurrensrätten gemensam , och inte att åternationalisera den .
Frågan om den enhetliga tillämpningen : vi skall vara medvetna om risken för en icke enhetlig tillämpning av konkurrensreglerna , men jag tror samtidigt att den risken inte skall överdrivas .
I likhet med flera andra föreskrifter i fördraget , artikel 81.1 och 82 , tillämpas de trots allt sedan decennier av nationella myndigheter och domare , och jag tycker inte att detta har skapat några större problem .
Inom ett överreglerat område är en enhetlig tillämpning i första hand beroende av graden av klarhet i de grundläggande rättsreglerna .
Kommissionen kommer att anstränga sig för att verkligen precisera den rättsliga ramen , såväl via allmänna åtgärder som i de praktiska besluten .
För det andra måste vi få till stånd effektiva konfliktförebyggande mekanismer och här föreslås i vitboken system för information och samråd .
Låt mig i det sammanhanget säga ett ord om den i mitt tycke utmärkta idé som framförts av Riis-Jørgensen och Huhne , dvs. idén om tillämpningsövervakning - monitoring of the implementation .
Så detta är vad idén att övervaka verkställandet går ut på .
Jag måste säga att jag tycker att det är en mycket god idé som vi troligen kommer att ta upp .
Även om vi har stor respekt för de nationella konkurrensmyndigheternas arbete och så vidare är det uppenbart att vi kommer att syna hur EG : s lagar tillämpas av nationella myndigheter och domstolar mycket noggrant .
Det är därför kommissionen vill ha kvar rätten att dra tillbaka ett fall från en nationell konkurrensmyndighet vid eventuell felaktig tillämpning .
Detta borde minska er oro i någon mån , fru Peijs .
( EN ) Vad beträffar Evans fråga om konsekvenserna för företagen är det viktigt att den samhällsekonomiska kostnads-intäktsanalysen genomförs på ett seriöst sätt .
Syftet med att ge ut en vitbok är när allt kommer omkring att inhämta synpunkter från företag lika väl som från andra källor .
Vi har fått in många utmärkta påpekanden och bidrag som ger oss underlag för att göra en kostnads-nytto-analys för industrin .
Vi kommer att gå igenom allt detta material noggrant innan vi lägger fram ett förslag till ny lagstiftning .
Det finns en aspekt av konsekvenserna för företagen som är mycket viktig .
Denna togs upp av Thyssen , Peijs och Palacio Vallelersundi : frågan om små och medelstora företag .
Många talare har betonat detta .
Kommissionen är särskilt uppmärksam på de små och medelstora företagens rättssäkerhet .
Vi föreslår ett system som stärker de små och medelstora företagens rättssäkerhet betydligt .
Varför ?
Är detta enbart en politisk gest ?
Nej .
I systemet föreslår vi att våra grundläggande regler ändras på ett sådant sätt att de flesta små och medelstora företag kommer att omfattas av generella undantag , såsom vad beträffar de vertikala begränsningarna .
De flesta små och medelstora företag har faktiskt en marknadsandel på mindre än 30 procent .
Vi har en de minimis-notis där vi förklarar att eftersom små och medelstora företag inte är involverade i marknadsdominans omfattas de normalt inte av det stränga förbudet i artikel 81.1 .
Vi arbetar på ytterligare generella dispenser och riktlinjer som alla kommer att ta hänsyn till de små och medelstora företagens speciella situation , och vår vitbok om modernisering kommer också att förbättra för de små och medelstora företagen genom att för det första den byråkrati det nuvarande anmälningssystemet ger upphov till försvinner och för det andra genom att artikel 81.3 blir direkt tillämplig , vilket kommer att gynna speciellt de små och medelstora företagen .
( IT ) Den fjärde frågan gäller rättssäkerheten .
Naturligtvis , Evans , är rättssäkerheten - jag är den förste att hålla med om det - viktig för företagen , inte bara för juristerna som även spelar en mycket viktig roll i det europeiska konstruktionsarbetet .
Rättssäkerheten är viktig för företagen : detta är en fråga som ordföranden för utskottet för rättsliga frågor och den inre marknaden , Palacio Vallelersundi som jag vill tacka för att hon alltid behandlar frågorna som rör den inre marknaden på ett uttömmande vis , dvs. i detta fallet inklusive konkurrensfrågan - även i sitt senaste inlägg underströk betydelsen av .
Jag är övertygad om att detta förslag kommer att öka företagens rättssäkerhet , och detta av tre anledningar : det gör det möjligt att utan ett föregående beslut godkänna samtliga konkurrensbegränsande avtal som uppfyller villkoren om utvidgning , tack vare den direkta effekten av artikel 81.3 ; det skapar möjligheter att hjälpa företagen om det uppkommer tolkningsproblem , genom publicering av motiverade beslut ; det kommer att åtföljas av undantagsbestämmelser och riktlinjer i avsikt att förtydliga reglerna och garantera deras säkerhet .
( FR ) Thyssen nämnde också frågan om företagsjuristernas legala privilegium .
Låt mig endast erinra om att EG-domstolen avgjorde den frågan 1982 , det vet ni bättre än jag .
Denna rättspraxis är fortfarande giltig och det finns ingenting som gör det motiverat att ifrågasätta den .
Enligt vitboken skall frågan åter granskas med avseende på en aspekt : utbyte av sekretessbelagd information .
Vilka garantier företagen bör få är för närvarande föremål för diskussioner .
( IT ) Herr talman !
Jag kommer så till Rapkays betänkande och jag vill först tacka ledamot Rapkay för kvaliteten i arbetet och för det stöd som ges kommissionens 28 : e årsrapport om konkurrenspolitiken .
Jag tycker mig finna en betydande samsyn , men i Rapkaybetänkandet understryks vissa saker som det är vår skyldighet att beakta mycket noga .
Jag vill av tidsskäl här endast peka på två : den ena gäller en ytterligare ökning av öppenheten .
Detta parlament vet att vi alla anser att öppenheten är en mycket viktig fråga inom konkurrenspolitiken , och jag personligen har från första början hävdat detta , alltsedan den 1 september , dvs. den första dagen av min utfrågning inför utskottet för ekonomi och valutafrågor .
När det gäller konkurrenspolitikens internationella dimension kan jag bekräfta för er , ledamot Rapkay , att kommissionen är beredd att lägga fram en rapport i frågan för parlamentet , denna fråga som även Randzio-Plath har pekat på och inom ramen för vilken jag kan nämna att vi har upprättat mycket tillfredsställande bilaterala kontakter med motsvarande myndigheter i USA , Kanada , Japan och vi kommer att arbeta för att Världshandelsorganisationen skall anta konkreta regler på konkurrensområdet .
Jag vill lika varmt tacka er , ledamot Jonckheer , för ert betänkande om sjunde översikten över statligt stöd i Europeiska unionen inom tillverkningsindustrin och vissa andra sektorer .
Jag tänker inte här gå in på frågan om medbeslutande , men det beror inte på att jag inte anser den viktig .
Den frågan har en institutionell betydelse som naturligtvis går utöver frågan om konkurrensen .
Jag har med andra ord inte rätt att uttala mig i en fråga som naturligt hör hemma inom ramen för regeringskonferensen .
När det gäller era förslag , ledamot Jonckheer , så vet ni redan att mina avdelningar - även om det sker med de alldeles för små , men mycket kvalificerade personalresurser de förfogar över - arbetar aktivt med att ta fram ett register över de statliga stöden och ett poängsystem över statliga stöd .
Jag väntar också med spänning på resultatet av den åttonde översikten , som har följande etapper : den sammanställs av tjänstemännen nu , i januari , och antagande av kommissionen i mars 2000 , för att se om de senaste tendenserna bekräftas .
Jonckheer , Thyssen och Gemelli har nämnt kandidatländernas förberedelser inom området konkurrens och när det gäller de statliga stöden .
Låt mig bara helt kort säga att vi arbetar med dem mycket aktivt och konkret : kandidatländerna förbereder sig , de har redan infört samtliga lagar på konkurrensområdet och de håller på att inrätta respektive myndigheter .
Jag kan också nämna , när det gäller oron - som jag , som ni vet , delar - för energin och framför allt miljön , att vi håller på att avsluta arbetet med att revidera lagstiftningen när det gäller statligt stöd på miljöområdet .
Jag vill också understryka , när det gäller problemen med statliga stöd , den punkt som togs upp av bland andra Riis-Jørgensen , om ersättning för juridisk hjälp .
I april 1999 antog kommissionen en ny förordning om specifika regler för sådan ersättning .
Ni kommer snart att märka - detta kan jag garantera er - att vi verkligen kommer att tillämpa de reglerna .
Slutligen , herr talman , ett par ord för att varmt tacka ledamot Langen för hans betänkande , som är mer sektorsinriktat , men som är lika viktigt för diskussionen .
Jag kan säga att kommissionens rapport i frågan om de statliga stöden till metallindustrin , som bekant , inte omfattar de individuella beslut som fattats när det gäller undantagsförfarandet , som anges i artikel 95 i fördraget om Europeiska kol- och stålgemenskapen , eftersom det rör sig om beslut som hamnar utanför tillämpningsområdet för lagen om stöd till stålindustrin .
När det gäller de kommande åtgärderna avseende stödåtgärder inom järn- och stålindustrin , som träder i kraft från och med juli 2002 , kommer vi att kräva att man fortsätter tillämpa stränga regler , vilket är ett behov som även branschen själv verkar instämma i .
När vi har lagt fram vårt förslag i frågan om nya regler och när vi har valt den juridiska form som är lämpligast , så skall det bli mig en glädje att få presentera vår vision för er .
Och det , herr talman , som jag tar med mig hem efter denna debatt , en debatt som jag vill tacka parlamentet för , är ett förbehållslöst intellektuellt och politiskt stöd från Europaparlamentets sida för en konkurrenspolitik , en grundläggande uppskattning för det arbete som kommissionen utför och ett förtroende för att det arbetet kan fortsätta i framtiden , saker som jag är särskilt tacksam för .
Vi kommer att fortsätta , framför allt med utskottet för ekonomi och valutafrågor , men även generellt sett med parlamentet , att föra den interinstitutionella dialog som har inletts .
I det sammanhanget gladde mig er kommentar , Palacio : vi måste alla ro , och helst i samma riktning .
Konkurrensen är inte ett mål , som mycket riktigt Rapkay har påpekat , utan ett mycket viktigt instrument i vårt europeiska konstruktionsarbete .
Som von Wogau sade i början på debatten , är konkurrensen trots allt inte något abstrakt : den ligger i medborgarnas intresse , den utgör en grund för den sociala marknadsekonomin .
Låt mig också tillägga att i det europeiska konstruktionsarbetet har konkurrensen haft , och kommer att fortsätta att ha , ett samhällsvärde och inte bara ett ekonomiskt värde .
Tack , kommissionär Monti .
Jag förklarar den gemensamma debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Straffrättsliga bestämmelser till skydd för unionens ekonomiska intressen Nästa punkt på föredragningslistan är betänkande ( A5-0002 / 2000 ) av Theato för budgetkontrollutskottet innehållande parlamentets rekommendationer till kommissionen om inrättande av straffrättsliga bestämmelser till skydd för unionens ekonomiska intressen .
Herr talman !
År efter år har vi förstått , framför allt av Europeiska revisionsrättens rapport , att pengar ur Europeiska unionens budget går förlorade på grund av slöseri , dålig förvaltning , oriktigheter och rent av verkliga bedrägerier .
Dessa missförhållanden har parlamentet pekat på både länge och väl för att sätta i gång åtgärder som skall tjäna till att skydda de europeiska skattebetalarnas pengar , som unionens budget när allt kommer omkring livnär sig av .
Särskild uppmärksamhet ägnas där kampen för att klara upp , beivra och förhindra bedrägerier .
Skapandet av UCLAF via Task Force , fram till inrättandet av Byrån för bedrägeribekämpning ( OLAF ) var viktiga steg , liksom förordningen för att skydda gemenskapens ekonomiska intressen och de lokala kontrollerna .
Påföljder för de fall som upptäcks kan av unionen utdömas enbart inom det administrativa området .
Kommissionens återkrav av orättmätigt erhållna belopp har hittills bara rönt måttlig framgång .
Straffrättsliga åtgärder ligger inom medlemsstaternas behörighetsområden .
Eftersom de båda rättsliga aspekterna ofta överlappar varandra och åsidosättande av unionens budget tilltar på ett gränsöverskridande sätt , och även begås av den organiserade brottsligheten , är behörigheten oklar bland medlemsstaterna .
Härtill kommer skillnader i de enskilda nationella rättsbestämmelserna , liksom utdragna och rent av ouppfyllda ömsesidiga framställningar om rättshjälp .
Detta har inte heller den av Europeiska rådet 1995 undertecknade konventionen om straffrättsligt skydd för gemenskapens ekonomiska intressen och de båda följande protokollen ändrat någonting på .
För att träda i kraft måste den ratificeras av alla 15 medlemsstaterna .
Efter fem år har hittills bara fyra medlemsstater gjort det .
Detta stillestånd , som hotar att undergräva unionens trovärdighet , har förmått parlamentet att ge impuls till en europeisk åklagarmyndighet .
Därigenom skall det inte på något sätt skapas gränsöverskridande straffrätts- eller rättsordning .
Målet är snarare att utrusta unionen med specifika instrument för att skydda dess ekonomiska intressen , och detta under iakttagande av subsidiariteten .
Med dagens betänkande återupplivar vi denna tanke och riktar en uppmaning till kommissionen att lägga fram lagstiftningsförslag för att förverkliga detta mål .
Därvid kommer begäran från utskottet för rättsliga frågor och den inre marknaden i dess yttrande , samt begäran från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor att tas med .
Vi uttalar två rekommendationer , som härrör från skapandet av OLAF och skall säkerställa dess operativa och rättsliga effektivitet , öppenhet samt skyddet av individens rättigheter .
Till detta behöver vi - det är den första rekommendationen - en rättsakt , där åtalspunkter som skadar unionens ekonomiska intressen är registrerade och där de ledande principerna är förankrade .
I ett ändringsförslag förespråkar jag en tidsfrist fram till den 30 september innan kommissionen skall lägga fram sitt förslag .
Den andra rekommendationen gäller straff- och straffrättsliga förfarandet .
Kommissionen bör fram till den 31 maj 2000 - även detta ändrat av mig - föreslå en rättsakt om skapandet av en oberoende organism , som institutionellt är bunden till kommissionen , för att samordna och kontrollera OLAF : s vederbörliga undersökningsverksamhet .
Den redan existerande övervakningskommittén kan bara kontrollera oberoendet för direktören i ämbetet .
Förslaget till en sådan rättsakt bör innehålla en oberoende stadga för denna organism och definiera dess uppgifter , som begränsas till OLAF : s interna utredningar och laga åtgärder som rör Europeiska gemenskapernas ekonomiska intressen , samt dess förbindelser med de nationella myndigheterna .
Något inflytande på rättsskipningen i medlemsstaterna är fortfarande uteslutet .
Övervakningen av rättsakternas rättmätighet skall tas över av EG-domstolen .
Dessutom uppmanar vi den kommande regeringskonferensen att ta upp en debatt om att skapa en europeisk åklagarmyndighet för att skydda unionens ekonomiska intressen , om möjligt på grundval av den undersökning som gjorts av namnkunniga forskare och nu erkänts i huvudsak , den s.k. corpus juris , liksom de senare publicerade genomförbarhetsstudierna .
Ytterligare rekommendationer för detta projekt återfinns också i den andra rapporten från de vises kommitté .
Kommissionen , Barnier och Vitorino , liksom vissa medlemsstater , är också öppna för idén .
Jag ber er , kära kolleger , att rösta ja till detta betänkande , som budgetkontrollutskottet har antagit med stor majoritet .
Vi kan här återigen ge ett tecken till att parlamentet är aktivt för att förebygga misshushållning och i synnerhet bedrägerier , och bestraffa detta , där så krävs .
( Applåder ) Herr talman !
Jag är glad över att få ta del i debatten om detta betänkande och vill framföra mina gratulationer till Theato .
Jag anser att detta är ett betänkande , där samarbetet mellan utskotten har fungerat väl , och det resultat som vi i dag har fått ta del av , är ett nyktert och sansat betänkande om en synnerligen känslig fråga .
Ett nyktert och sansat angreppssätt är särskilt nödvändigt vad beträffar artikel 280.4 .
För om vi ville ge ett pris åt den artikel som är mest svårbegriplig , otydlig och oklar - eller vad man nu vill kalla det - så skulle konkurrensen garanterat vara mycket jämn , för fördraget består av en brokig samling komplicerade artiklar , men denna är utan tvekan en av de starkaste kandidaterna till ett sådant pris .
Samtidigt är det en synnerligen känslig fråga , eftersom det handlar om skyddet av gemenskapens ekonomiska intressen , så som Theato så riktigt uttrycker det .
Vi är alla medvetna om behovet - och parlamentet har tagit upp eller fört fram det problemet - av att skydda gemenskapens ekonomiska intressen .
Men se upp , som fransmännen säger , " ne jettons pas le bébé avec l ' eau du bain " , det vill säga , i skyddet av gemenskapens ekonomiska intressen måste man å ena sidan respektera - och det påpekar Theato - de nationella staternas behörighet , men även andra saker som påverkar medborgarna , sådant som påverkar de grundläggande garantierna .
Slutsatserna i Theatos betänkande värnar om dessa .
Därför hoppas jag i egenskap av ordförande för utskottet för rättsliga frågor och den inre marknaden , och givetvis även som ledamot , att parlamentet i morgon antar betänkandet med stor majoritet och att kommissionen verkställer det på bästa sätt .
Herr talman !
Som Theato sade är detta ett kritiskt betänkande .
Det är ett betänkande som har föreslagits av budgetkontrollutskottet och det är ett initiativbetänkande .
En av anledningarna till att vi var mycket angelägna om att lägga fram detta var att Europeiska unionen , vare sig vi tycker om det eller inte , är beryktad för bedrägerier och misskötsel .
Detta är ibland överdrivet men så är det .
Vi måste göra någonting åt det .
En del av medlemsstaterna har inte åtföljt vissa av de åtgärder vi har vidtagit tidigare - och låt oss inte glömma att medlemsstaterna svarar för verkställandet av omkring 80 procent av EU-budgeten .
Många av dem har inte undertecknat , eller inte ratificerat konventionen om skyddet av ekonomiska intressen , och därför stod det klart att något mer radikalt behövde göras .
Vi måste ta detta ansvar på allvar .
Vi måste kunna åtala människor som begår bedrägerier gentemot Europeiska unionen .
Frågan är : vem skall åtala ?
Det är här vi verkligen kommer i problem .
Vems ansvar är det när det rör sig om ett organ som överskrider så många gränser ?
Vi måste också ta hänsyn till medlemsstaternas oro .
Förslaget att etablera en europeisk allmän åklagarmyndighet är mycket känsligt .
Vi är alla medvetna om att en helhjärtad federalistisk inställning och en situation där en europeisk juridisk myndighet står över de nationella juridiska myndigheterna enligt vissa är att gå för långt .
Men diskussionen måste starta och vi uppmanar därför regeringskonferensen att inleda diskussioner .
Det viktigaste för parlamentet , i egenskap av Europeiska unionens budgetövervakare , är hur man skall handskas med anställda inom Europeiska unionens institutioner .
I en tid då vi ser över hela reformprocessen är det avgörande att vi ger rätt signaler .
Människor måste inse att om de begår bedrägerier kommer de att åtalas , så är inte fallet för närvarande .
Hela frågan om vi har laglig befogenhet att göra detta har Palacio skisserat .
Jag skulle vilja slå fast att min grupp kommer att föreslå en ändring som innebär att passusen om hur kommissionen bör handskas med denna fråga tas bort .
Vi är medvetna om att detta är en känslig debatt .
Vi vet att kommissionen kanske behöver spelrum för att förhandla fram en situation som alla parter kan acceptera .
Låt mig bara göra klart att vi inte förbinder oss till en corpus juris här , inte förbinder oss till en europeisk allmän federal åklagare .
Men vi förbinder oss definitivt att förändra ett status quo som är helt oacceptabelt .
Herr talman !
Jag skulle vilja börja med att lyckönska fru Theato till hennes betänkande .
Jag anser att det är ett utmärkt betänkande och att den övervägande delen av det kommer att stödjas av min grupp .
Men jag får en stark känsla av att hon på detta stadium egentligen hade velat gå ett steg längre .
När jag lyssnat till diskussionerna under de senaste fem , sex månaderna skulle det mycket väl kunna vara fallet .
Vi vet alla att vi 1995 kom överens om att man måste sörja för ett bättre straffrättsligt skydd för unionens ekonomiska intressen .
Men medlemsstaterna var inte med på noterna .
Det är helt enkelt ett politiskt faktum , och enligt vad jag tror kan vi för närvarande inte göra mycket åt detta .
Den möjlighet som nu finns är att kommissionen på grundval av artikel 280 i fördraget tar nya initiativ , och jag skulle vilja föreslå kommissionen att verkligen göra detta så snabbt som möjligt .
Min grupp är , i motsats till föregående talare som redan försvunnit , en stark förespråkare för en europeisk allmän åklagare .
Min kollega Jan-Kees Wiebenga kommer utan tvivel att ytterligare gå in på detta , för han har tidigare författat ett betänkande i ämnet .
Det som vi har behov av , tror jag , är en definition på europeisk nivå av vad som exakt menas med bedrägeri och oegentlighet .
Jag var själv med i undersökningskommittén om transittrafiken .
Ett av de stora problemen på det området var att om man gör något fel , och då handlar det framför allt om Europeiska unionens inkomster , så är det en oegentlighet i det ena landet och ett brott i det andra landet .
Så kan vi inte ha det längre tyckte jag , i synnerhet inte för närvarande .
En allmän politisk punkt .
Något som vi också kan konstatera i fråga om Europavalet är att det låga valdeltagandet är ett faktum .
Vi kan förbättra detta genom att snabbt ta itu med brottsligheten i Europa , och det måste ske på europeisk nivå .
Herr talman !
Även mitt tack går till föredraganden .
Theatos betänkande kan bidra till att det åter skapas förtroende för de europeiska institutionerna .
Jag tror att vi alla verkligen behöver det , om vi tänker på resultaten från de senaste Europavalen , och på valdeltagandet .
Det är ju samma problem varje år .
Revisionsrätten offentliggör sin rapport , och i rapporten beskylls medlemsstaterna för olika bedrägerier .
Men de europeiska institutionerna har hittills haft alltför få möjligheter att ingripa och se till att något verkligen görs , att det avhjälps .
Just detta förfarande minskar förtroendet varje år på nytt .
Jag tror att Theatos betänkande och hennes förslag kan bidra till att situationen vänder , och att det klargörs att de europeiska institutionerna ser till att de europeiska pengarna också satsas målinriktat och att det här inte förekommer några bedrägerier .
Det är viktigt att vi efter det första steget som redan tagits , nämligen att ur UCLAF skapa OLAF , en oberoende institution , nu tar ett andra steg och även skapar en rättslig ram för OLAF , så att OLAF kan agera inom en säker rättslig ram .
Till detta behöver vi den europeiska åklagarmyndigheten , som ser till att det finns en klar rättslig garanti , även för de misstänkta .
Jag måste dock säga att min grupp tyvärr inte kommer att rösta enhälligt för ert betänkande .
Jag hoppas att debatten kommer att övertyga ytterligare några personer .
Betänkligheterna är tyvärr fortfarande alltför stora för att det här kommer att skapas en europeisk institution , som minskar subsidiariteten .
Men jag vill bidra med min del så att Theatos betänkande skall få ett större stöd .
Herr talman !
Vi är i allt väsentligt positiva till den resolution som lagts fram även om vi anser att detta inte kan bli annat än en uppmaning från parlamentet till rådet att genom en ändring av fördragen se till att skapa ett effektivt straffrättsligt skydd för unionens ekonomiska intressen .
Inrättandet av en europeisk åklagare och tillskapandet av brottsrubriker som är gemensamma för samtliga länder inom unionen är utan tvekan en god idé , men jag anser det vara omöjligt att försöka förverkliga den utan att först ha inrättat en gemensam rättsordning för unionen .
Vi talar ju här om straffrätten , det område där motståndet från nationalstaterna mot gemensamma regler är och alltid har varit starkt .
Det är i själva verket otänkbart att man skulle kunna skapa gemensamma straffrättsliga regler för en enda sektor , nämligen skyddet av ekonomiska intressen , utan att först ha skapat ett gemensamt europeiskt rättssystem .
Det räcker att man läser de exakta och uttömmande motiven i Theatos betänkande för att man skall inse vilka problem som återstår att lösa .
Men idén bör uppmuntras och det råder ingen tvekan om att man under dessa försök att skydda de ekonomiska intressena upptäcker behovet av att inrätta en gemensam corpus juris och att införa den i fördragen .
För egen del och som företrädare för min grupp vill jag också framföra en förhoppning om att unionens ekonomiska intressen blir en vägröjare för insikten om att det behövs ett europeiskt rättssystem som respekterar medborgarnas garanterade rättigheter , dvs. ett rättssystem som lyfter fram de garantier som , dessvärre , i många medlemsstater inte har nått upp till en godtagbar nivå .
Jag uttrycker därför , som företrädare för min grupp , min uppskattning av Theatos betänkande .
Men jag anser att det i grunden handlar om en fråga som måste föras upp på dagordningen för regeringskonferensen .
Herr talman !
I betänkandet av Theato om skyddet av Europeiska unionens ekonomiska intressen föreslås bl.a. att man , i första hand , skall centralisera de straffrättsliga processerna genom att inrätta en europeisk åklagarmyndighet .
Detta förslag står helt uppenbart i strid med andan i det nuvarande systemet , där straffrätten och straffrättsliga processer - centrala element i de nationella rättssystemen - skall lyda under varje folks suveränitet och varje stats exklusiva ansvarsområde .
Idén om en europeisk åklagarmyndighet syftar tvärtom till att på sikt begränsa staterna och ge dem en underordnad roll i de här frågorna .
Dessutom skulle förslaget utlösa en räcka reformer som är helt omöjlig att förutse .
Enligt Theatobetänkandet skulle en europeisk åklagarmyndighet vara nödvändig , bl.a. för att förbättra ledningen av undersökningarna vid Byrån för bedrägeribekämpning , OLAF .
Men samtidigt får vi veta , i betänkandet av Van Hulten som diskuteras i dag , att den europeiska åklagarmyndigheten själv skall övervakas av en domstol i Europeiska unionen .
På så sätt kan en liten europeisk reform dölja en medelstor , och en medelstor dölja en stor .
Och då räknar jag inte med att en stor reform i sin tur kan dölja en gigantisk reform , eftersom vi snart kommer att få se ett förslag till en europeisk straffrätt och varför inte - på sikt - en europeisk justitieminister som kontrolleras genom en utvidgning av Europaparlamentets befogenheter .
Jag tror således att vi borde reflektera över den maktbalans som man riskerar att kullkasta genom att presentera reformer av det här slaget , vilka kan framstå som avgränsade .
Slutligen anser vi att den här typen av förslag , såsom förslaget om en europeisk åklagarmyndighet , avslöjar en oförmåga att föreställa sig Europa på något annat sätt än i en pyramidisk och centraliserad form , organiserad kring en överstat .
Gruppen Nationernas Europa vill tvärtom ha ett Europa med många centra som binder samman nationerna i ett nätverk .
Detta nät skulle t.ex. kunna innebära en bättre samordning mellan nationella åklagarmyndigheter , och man skulle eventuellt kunna inrätta nationella utbildningar med inriktning på brott som skadar gemenskapens finanser .
Herr talman !
Det finns således redan en juridisk struktur , och dess principer är bra .
Vi behöver endast fullända den .
Herr talman !
Theato föreslår en institutionell revolution av två skäl .
Allmänheten påstås vara likgiltig inför 20 miljoner arbetslösa och tusentals galna kor , men oroad över de bedrägerier som äventyrar de ekonomiska intressena , och dessa två skäl skulle motivera två bestämmelser : en europeisk straffrätt om anti-gemenskapliga förbrytelser och en europeisk allmän åklagarmyndighet .
Theato har förresten , sannolikt , glömt ett europeiskt fängelse , eftersom FBI - den europeiska polisen - existerar i och med OLAF .
Allt detta skulle inrättas genom två förordningar , en för åklagarmyndigheten och en för straffrätten .
Det är förordningar som antas på grundval av artikel 280 i fördraget , dvs. med utgångspunkt i den avledda rätten , för det som utmärker den avledda rätten är att man tillåter alla strömningar som leder i andra banor .
Det finns faktiskt två strömningar .
Först och främst den klassiska ideologiska , eurofederalistiska strömningen : för en gemensam marknad , en gemensam mervärdesskattesats , en gemensam diplomati , en gemensam armé och nu en gemensam straffrätt och en gemensam åklagare .
Allt detta för att bekämpa bedrägerier som underskrider en miljard euro , samtidigt som man mister tiotals miljarder euro på grund av allmänna preferenssystemet , frihandelsområdena , tullgåvor till Chiquita och miljarder som förlorats på den fjärde resursen , BNI , ett resultat av pakten om finansiell åtstramning .
Sedan har vi den puritanska strömningen ; det nordtyska Europa , det lutheranska och calvinistiska Europa , Kväkareuropa , som vill påtvinga oss sin moraliska ordning .
För i grunden är det så , att ju mer man lättar på seder och bruk , desto hårdare håller man i plånboken .
Herr talman , mina damer och herrar !
Det är absolut nödvändigt med ett verksamt straffrättsligt skydd för Europeiska unionens intressen , i dag mer än någonsin .
Bedrägeri- och korruptionsskandalerna i det förflutna har på lång sikt skakat förtroendet hos Europas medborgare .
Trovärdigheten i de ansträngningar vi gör här i parlamentet för att de ekonomiska medlen skall satsas korrekt står och faller med våra ansträngningar för att behandla dem och förhindra dem i framtiden .
Hit hör inte bara administrativa , utan också strukturella förändringar , dvs. vi måste skapa de instrument med vilka man över huvud taget kan garantera ett straffrättsligt skydd .
Regeringskonferensen 2000 är lämplig som diskussionsforum för detta .
Nu kan man naturligtvis inta den ståndpunkten att straff- och straffprocessrätten hör till medlemsstaternas rättssystem och inte kan röras när man har en subsidiaritetsprincip .
Själv hör jag utan tvivel till dem som förfäktar denna princip och till motståndarna av all vidare utvidgning av de europeiska ansvarsområdena .
Just i samband med kraven på regeringskonferensens arbete bör tyngdpunkten ligga på att fordra en klar ansvarsavgränsning .
Men detta innebär inte någon motsägelse , ty när man kräver ett straff- och straffprocessrättsligt instrument , så som anförs i betänkandets rekommendation I och II , handlar det egentligen om att iaktta EU : s ursprungliga egna intressen , som såtillvida inte skadar medlemsstaternas rättsliga intressen , utan tvärtom stöder dem , åtminstone indirekt .
Förenligheten med de olika nationella rättssystemen , som bekräftats av experterna , visar att man i Europa har mycket gemensamt även på det straffrättsliga området , exempelvis när det handlar om innehållet i de här tillämpliga åtalspunkterna .
Med hänsyn till dessa synpunkter anser jag att skapandet av en sådan ram som krävts är riktigt och också är påbjudet som en vidareutveckling av OLAF .
Herr talman !
Kommer en europeisk offentlig åklagare att kunna avskaffa fotbollsbedrägerierna med EU-medel ?
Jag tror inte det .
Vi kan istället komma långt med de befintliga instrumenten .
Eurojust skulle kunna vara ett alternativ till den europeiska offentliga åklagaren , vilket föreslogs på det senaste toppmötet .
Eurojust skall i inledningsskedet lyda under Europol och stödja forskningen i brottsfrågor .
Det är precis ett sådant praktiskt samarbete det finns behov av .
OLAF , Europol och konventionen om utlämning och ömsesidig rättshjälp skall utnyttjas fullt ut , och när bedrägerikonventionen från 1995 slutligen blir ratificerad av medlemsstaterna , kan vi även komma långt med hjälp av den .
Jag håller emellertid med föredraganden : Det är fullständigt oacceptabelt att de flesta medlemsstaterna ännu inte har ratificerat den .
Det är helt enkelt för dåligt och jag förstår mycket väl att folk blir otåliga och kräver att vi i stället skall få en gemensam europeisk åklagare .
Det är emellertid en stor mastodont att bygga upp .
Det är ändå bara de grövsta fallen som kommer att få straffrättsliga konsekvenser .
90 procent av fallen kommer att utgöra disciplinfrågor om försummelse eller inkompetens .
I stället finns det behov av en ordentlig intern kontroll och bättre möjligheter att avskeda folk .
Vi skall ändra tjänsteföreskrifterna och det disciplinära förfarandet och inte minst skall vi ändra praxis .
För närvarande används aldrig artikel 52 i tjänsteföreskrifterna om avskedande på grund av grov försummelse .
Skall vi inte se till att rensa upp ordentligt och hålla rent framför vår egen dörr , innan vi förhastar oss och börjar bygga upp nya förkromade institutioner ?
Herr talman !
Vi vill allesammans gärna göra något för den europeiska bedrägeribekämpningen .
Men frågan är nu : gör Europeiska unionen också något för denna ?
Svaret är att vi vet alldeles för litet om detta .
Toppmötet i Tammerfors handlade om brottsbekämpning .
Alla var så kallat nöjda med detta , men i själva verket gjordes det inte några större framsteg .
Det finns fortfarande ingen gällande europeisk antibedrägerilagstiftning , eftersom medlemsstaterna , vilket redan har sagts , inte har ratificerat de framlagda fördragstexterna .
På det området måste det således hända mycket .
Och vad är det då som måste hända ?
Det är två saker , och i Theatos betänkande framkommer detta på ett klart och tydligt sätt .
För det första , i alla Europeiska unionens medlemsstater måste samma straffbestämmelser gälla i fråga om europeiskt bedrägeri .
Likriktning på detta begränsade område .
För det andra måste verkligen en europeisk åklagarmyndighet inrättas , och den skall ha två uppgifter : för det första att stödja de nationella allmänna åklagarna , att hjälpa till med åtal i fråga om europeiska bedrägerimål , och för det andra att övervaka Europol och OLAF i rättsligt avseende , för detta är två utredande myndigheter som för närvarande kan operera okontrollerat i rättsligt avseende .
Den europeiska åklagarmyndigheten är inte någonting att vara rädd för ; det jag hör här runt omkring mig är bara skräckscenarior .
Det är helt enkelt något mycket positivt , precis som Europol .
Europol , polissamarbetet , står inte över de nationella polismyndigheterna , utan finns med tanke på informationsutbytet mellan polismyndigheterna .
Det är precis på det sättet som en liten begränsad europeisk åklagarmyndighet måste börja arbeta .
Det gäller inte bara under uppspårningsfasen , utan också under åtalsfasen .
Parlamentet är för detta .
Den oberoende expertkommittén är för detta .
Jag uppmanar ministerrådet och Europeiska kommissionen att också erkänna denna åtgärd .
Herr talman !
Jag skall koncentrera mig på frågan om corpus juris .
Jag vill verkligen stödja det Morgan sade om detta .
Corpus juris är någonting som sattes ihop utan någon offentlig debatt eller deltagande alls .
Tanken med en europeisk allmän åklagare med överordnad jurisdiktion inom EU : s territorium skulle få stora konsekvenser för de traditionella systemen både i Irland och i Storbritannien .
Planerna på en enda strafflagstiftning och en europeisk allmän åklagare är någonting medlemsstaterna har rätt att få information om .
När planen först gjordes upp sade de att den skulle vara begränsad till fall av bedrägeri mot EU : s budget .
Men när corpus juris lanserades i San Sebastian 1977 - inför en mycket utvald publik på 140 jurister , utan inbjudna media - sade den dåvarande talmannen i Europaparlamentet , Gil-Robles Gil-Delgado , att han ansåg att den var på embryostadiet och att avsikten var att utvidga EU : s befogenheter på brottsmålssidan till att omfatta all kriminell verksamhet .
Vi behöver en offentlig debatt om detta .
Medlemsstaterna och medborgarna i medlemsstaterna måste få ordentlig information .
Frågan om hotet mot det traditionella juridiska systemet i Irland och Storbritannien måste tas upp .
Det behövs mycket större öppenhet och insyn än hittills i denna fråga .
Det är oacceptabelt att någonting dylikt har prackats på EU : s medlemsstater utan någon ordentlig offentlig debatt .
Herr talman , kära kolleger !
I budgetkontrollutskottet avstod jag från att rösta om denna text i min egenskap av företrädare för de radikala ledamöterna , för jag delar den oro som på ett så kunnigt vis formulerats av företrädaren för en annan mycket viktig juridisk tradition , dvs. den som har formen av common law .
Med den här texten rör vi oss verkligen i utkanten av vad som är möjligt , eftersom vi anser att det finns frågor som måste lösas och att det är viktigt att bedrägerierna inom gemenskapen stoppas , att de stryps .
Men det sätt på vilket vårt utskott , tack vare ordföranden Theatos energi och envishet , har för avsikt att förverkliga intentionerna i denna text får inte ske utan kritik .
En annan viktig kritik som kan riktas mot texten gäller sekundärrätten .
Artikel 280 i fördraget ger rådet rätt att bestämma om lämpliga instrument för att bekämpa bedrägeriet .
Men vi blir ändå en aning förvånade över att man vill inrätta en institution , vilket innebär ett kvalitetssprång , utan att genast kunna förutse vilka motåtgärder som kommer , dvs. man bortser från försvaret och därmed möjligheten att åklagare och försvarare skall kunna fungera effektivt i ett så viktigt rättssystem .
Genom att avstå från att rösta i utskottet har vi velat uttrycka denna vår tveksamhet .
Herr talman !
Jag tror att det är något som måste sägas tydligt i denna fråga i denna församling , i plenarsammanträde och i utskotten , eftersom det är uppenbart att debatten inte får bortse från den kulturella bakgrunden , den juridiska kulturen och de miljöer i vilka de institutionella frågorna skall tas upp .
Vi står inför mycket allvarliga händelser som i det förflutna verkade vara en tradition .
I dag har något förändrats , åtminstone när det gäller mekanismerna , framför allt när det gäller kontrollen , men vi är ändå inte nöjda , framför allt inte om man i berörda fora pratar om en europeisk åklagare , brott , bedrägerier , förskingring och avslöjanden av hemligheter på europeisk nivå .
Jag anser naturligtvis att vi måste skydda gemenskapens intressen och dess rykte , förutom relationerna med bidragsgivarna , som utgör en omistlig och avgörande del av gemenskapens liv .
Av den anledningen är det riktigt att undersöka frågan om ett skydd av intressen av mer allmän och universell natur , och att på ett bättre sätt förena sig med rättssystemen inom de enskilda staterna .
I det sammanhanget uppstår en känsligare fråga : hur förhåller sig en europeisk åklagare till de enskilda medlemsstaterna och det rättssystem som är uppbyggt inom ramen för dem ?
Detta är en fråga som fortfarande måste tas upp såväl ur kulturell som praktisk synpunkt .
I dag riskerar vi att lägga en ny institution ovanpå de många skilda institutioner som redan existerar i de enskilda länderna .
Herr talman !
Jag vill gärna helt snabbt säga något om två punkter .
För det första : Jag vill inte referera till de filosofiska frågorna om medlemsstaternas subsidiaritet och suveränitet , även om jag absolut anser att en sådan debatt bör föras , eftersom mitt regelbundna tittande på brittiska TV-sändare ändå får mig att inse vad nationella politiker där betraktar som ett hot mot den inhemska rättskulturen från kontinentens sida .
Ibland är det nästan kabarébetonat och förtjänar att diskuteras .
Men det är inte det jag vill tala om .
Jag vill tala om Theatos betänkande .
Jag tror att man har trasslat in sig i de juridiska svårigheter som finns här - och uppenbarligen finns det bara en mycket liten möjlighet för Europeiska unionen att ta upp dessa åtalspunkter som europeiska åtalspunkter .
Jag refererar till rekommendationerna 1 och 2 .
Det står ju där inte längre något om en europeisk åklagare , utan av juridiska orsaker har det nu blivit en oberoende europeisk myndighet , med Theatos ord tidigare en organism .
Där har vi uppenbarligen problem med den rättsliga grunden .
Sedan har vi problem med åtalspunkterna .
Det har inte ändrats .
Där finns det fortfarande åtalspunkter , som så att säga också går utöver de europeiska åtalspunkterna , eller åtminstone kan gå utöver dem , exempelvis penningtvätt , häleri och stämpling .
I det avseendet anser jag att det finns juridiska oklarheter , som bör undanröjas .
Men det som är absolut nödvändigt , och därför kommer vi att rösta för punkt 1 utan dessa rekommendationer , är en klar politisk signal från parlamentet till kommissionen och rådet att vi med hjälp av en klar rättsakt vill ha ett slut på de förhållanden , som har gripit omkring sig .
Herr talman !
Parlamentet har sedan flera år krävt en specifik och enhetlig straffrätt till skydd för unionens ekonomiska intressen .
Sanningen är att frustrationen ökar när vi konstaterar svagheterna i konventionen ( och protokollen i anslutning till detta skydd ) , som fem år efter att den undertecknats ännu inte har ratificerats eller trätt i kraft .
Mer voluntaristiska försök , som det nuvarande OLAF , övervinner inte den legitima oron över garantisystemet för de individuella rättigheterna .
Förslagen i Theatos betänkande för att uppmuntra kommissionen att lägga fram en rättsakt om straffrättsliga bestämmelser till skydd för unionens ekonomiska intressen med typfall för brott , framför allt oredlighet avseende bidrag från och avgift till gemenskapens budget , är enligt vår mening ett försök att införa en ny och allt nödvändigare enhetlig straffrätt i gemenskapen .
Samtidigt är de en vädjan om inrättande av ett " oberoende europeiskt organ " , som samordnar och kontrollerar att OLAF : s utredningsverksamhet följer gällande bestämmelser , utan att det påverkar medlemsstaternas rättskipning och under EG-domstolens övervakning .
Slutligen , i Tammerforsbeslutens fotspår tas i betänkandet återigen ett europeisk åklagarämbete upp , vilket kommissionär António Vitorino i ett lämpligt ögonblick beslutade sätta ljuset på genom att begära att regeringskonferensen skulle ta upp skapandet av denna nya tjänst i sin dagordning , det ämbete som alla i dag anser är nödvändigt .
Eftersom behovet av rättslig och effektiv disciplin i institutionerna vidhålls , genom att tillsluta unionens ekonomiska system med en europeisk materiell och processuell rätt anpassad till förtroendet för gemenskapens ekonomiska liv , stöder vi detta betänkande .
Emellertid finns det några mycket enkla frågetecken .
Finns det tillräckligt med rättslig grund för att motivera skapandet av en ny specifik straffrätt för gemenskapen som , även om man kan kalla den subsidiär , i praktiken och i vissa områden alltid kommer att strida mot medlemsstaternas traditionella och partiella straffrätt ?
Skulle det inte vara mer politiskt korrekt , när det råder tvivel , att föra upp reformen av rättssystemet på regeringskonferensens dagordning , och alltså ta upp dessa förslag i den mer allmänna reformen av unionens rättssystem , och ta upp dem i den bild man vill ge den europeiska åklagaren ?
Är inte dessa frågor av största intresse för en revidering av fördragen som kan bidra till att befästa området med frihet , säkerhet och rättvisa i unionen ?
Herr talman !
EU utsätts i dag för hård granskning .
Förtroendet för unionen är allvarligt skadat .
För att råda bot på detta krävs krafttag .
Vi välkomnar därför ökade resurser till OLFAF , så att vi effektivare kan utreda alla misstankar .
Vi ser det samtidigt som självklart att de som begår brott mot EU på ett effektivt sätt måste kunna ställas till ansvar .
Det är beklagligt att konventionen om skydd för unionens ekonomiska intressen har genomförts i så få medlemsstater .
Vi menar därför att det är rimligt att kommissionen får i uppdrag att lägga fram förslag , som innebär att den rättsliga ram som redan finns vidareutvecklas .
Däremot är jag inte övertygad om att en sådan effektivisering kräver en gemensam europeisk lagstiftning eller en centralisering av sådan brottsbekämpning .
I dagsläget är jag därför skeptisk till idén om en europeisk åklagare , vilken knappast är möjlig att genomföra inom ramen för dagens fördrag .
Vi tror mer på Eurojust , där nationella åklagare samarbetar .
Det stora problemet är inte att brott mot unionen inte beivras , utan att de så ofta begås och alltför sällan upptäcks .
Utmaningen för kommissionen och för oss är dock att finna rätt mix .
De bedrägerier och den misshushållning som förekommer får inte leda till att vi fastnar i en ålderdomlig hierarkisk byråkrati , som genom överdriven detaljkontroll förhindrar utvecklingen av modern förvaltning .
Därför välkomnar vi den offensiva synen i Van Hultenbetänkandet .
Huvudlinjen bör vara att varje förvaltning tar ansvar för sin egen kontroll .
Våra erfarenheter av modern förvaltning säger oss att öppenhet , decentralisering av ansvaret och kvalificerad utvärdering ofta är lika effektivt som byråkratisk detaljkontroll .
Den stora utmaningen är därför att skapa en modern och effektiv förvaltning utan att förlora i rättssäkerhet och kontroll .
Det kräver personalutbildning , modernare rekryteringsmetoder och framför allt öppenhet och insyn .
Att kunna granska förvaltningen effektivt är det bästa skyddet mot oegentligheter .
Herr talman , fru föredragande , ärade ledamöter !
Att skapa nytt förtroende från medborgarnas sida för de europeiska institutionernas arbete och nytt förtroende för den europeiska politiken , är en av de viktigaste uppgifter vi står inför .
Kommissionen har åtagit sig denna uppgift , och utkastet till det totala paketet med de inre reformerna dokumenterar detta .
Parlamentet har åtagit sig denna uppgift , och föreliggande betänkande utgör ett imponerande bevis för det .
Jag vill ge föredraganden kommissionens erkännande för att hon på nytt har ägnat sig åt den verkligt svåra frågan om vilka rättsliga grunder , vilka institutionella ändringar som kan göras för att intensifiera bekämpningen av de bedrägerier som drabbar Europeiska unionen .
Alla medlemsstater har i och med ratificeringen av Amsterdamfördraget intygat att de vill ge bekämpningen av bedrägerier mot Europeiska unionens ekonomiska intressen samma prioritet som bekämpningen av bedrägerier som drabbar dem själva , men i realiteten har fortfarande enbart de första fyra medlemsstaterna ratificerat det 1995 beslutade avtalet .
Kommissionen är helt överens med föredraganden om att denna situation inte är acceptabel .
En rättsakt , ett direktiv , där åtalspunkter i samband med bedrägeri , exempelvis penningtvätt eller korruption , definieras enhetligt och där förpliktelsen till rättsliga åtgärder fastställs som ett bindande mål , kan här innebära ett viktigt steg , och jag kommer därför att föreslå kommissionen att den mycket snart skall granska detta steg .
OLAF , den europeiska byrån för bedrägeribekämpning , är ett av kommissionens viktigaste instrument för att uppfylla sitt åtagande att bekämpa bedrägerier .
Kommissionen har därför inte accepterat att de båda europeiska bankerna Europeiska centralbanken och Europeiska investeringsbanken har bestridit OLAF : s rätt att undersöka även dessa båda institutioner , under hänvisning till sin oberoende ställning .
Kommissionen har därför vid sitt senaste sammanträde beslutat om ett överklagande mot dessa båda banker , och jag hoppas att parlamentet godkänner denna åtgärd .
Den andra rekommendationen i föreliggande betänkande gäller granskningen av rättmätigheten i OLAF : s undersökningsåtgärder i de olika europeiska institutionerna .
Övervakningskommittén för OLAF , som inrättades samtidigt med OLAF , har till uppgift att säkerställa OLAF : s oberoende , men den kan inte utöva den verksamhet som nämns i betänkandet , att kontrollera OLAF : s interna utredningsarbete .
Här är jag fullständigt överens med övervakningskommittén och med föredraganden .
Det betyder att det här finns en brist som måste åtgärdas , och jag kommer med tanke på en vidareutveckling att granska den väg som föreslås i betänkandet .
Jag vill dock be om en sak : Jag tror att man måste förhindra att debatten om en utvidgning av den rättsliga grunden för OLAF leder till missuppfattningen att OLAF nu inte skulle ha tillräcklig auktoritet .
Nej , det får inte leda till att OLAF : s auktoritet undergrävs , och jag tror inte heller att föredraganden avser det .
Därför ber jag er att helt och fullt stödja OLAF : s arbete även i dess nuvarande form .
( Applåder ) Tack , kommissionär Schreyer .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
OMRÖSTNING ( Parlamentet godkände kommissionens förslag . )
Heaton-Harris ( PPE-DE ) .
( EN ) Herr talman !
Som en ordningsfråga skulle jag vilja be er om ett klargörande av arbetsordningen , nämligen artiklarna 133.2 och 138.4 .
De handlar båda om omröstning .
Är det inte så att vid andra omröstningar än omröstningar med namnupprop skall omröstning först ske genom handuppräckning och först sedan , om det finns tvivel om utgången , skall vi använda det elektroniska voteringssystemet ?
Kära kollega !
Det stämmer att jag genomförde en omröstning med handuppräckning , eftersom ingen grupp hade begärt en omröstning med namnupprop .
Som ni vet genomförs endast omröstningar med namnupprop och elektroniska omröstningar om kollegerna begär detta .
I det här fallet kan jag försäkra er att det fanns en överväldigande majoritet för det direktiv som vi just har röstat igenom .
Herr talman , jag syftade inte på just denna omröstning utan på omröstningar i allmänhet .
Det är uppenbart att vissa ordförande inte tittar på händerna , så att säga , utan går direkt till det elektroniska voteringssystemet .
Jag undrade om detta är ett korrekt tillvägagångssätt .
Jag vet att det tar längre tid , men borde vi inte alltid först räcka upp händerna ?
Jag försäkrar er , kära kollega , att jag kommer att vara mycket uppmärksam på hur många händer som räcks upp .
Jag hoppas att det blir många då det är dags för omröstning .
Förslag till Europaparlamentets och rådets direktiv om tillnärmning av medlemsstaternas lagstiftning om märkning och presentation av livsmedel samt reklam för livsmedel ( kodifierad version ) ( KOM ( 1999 ) 0113 - C4-0212 / 1999 - 1999 / 0090 ( COD ) ) ( Utskottet för rättsliga frågor och den inre marknaden ) ( Parlamentet godkände kommissionens förslag . )
Förslag till rådets förordning ( EG , Euratom ) om genomförande av beslut 94 / 728 / EG , Euratom om systemet för gemenskapernas egna medel ( kodifierad version ) ( KOM ( 1997 ) 0652 - C4-0018 / 98 - 1997 / 0352 ( CNS ) ) ( Utskottet för rättsliga frågor och den inre marknaden ) ( Parlamentet godkände kommissionens förslag . )
Förfarande utan debatt Betänkande ( A5-0106 / 1999 ) av Varela Suanzes-Carpegna för fiskeriutskottet om förslag till rådets förordning om slutande av det protokoll i vilket de fiskemöjligheter och finansiella motpartsmedel fastställs som föreskrivs i avtalet mellan Europeiska ekonomiska gemenskapen och Demokratiska republiken São Tomé och Príncipes regering om fiske utanför São Tomé perioden 1 juni 1999 - 31 maj 2002 ( KOM ( 1999 ) 0550 - C5-0305 / 1999 - 1999 / 0228 ( CNS ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Andrabehandlingsrekommendation ( A5-0105 / 1999 ) från utskottet för regionalpolitik , transport och turism om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets direktiv om harmonisering av examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg eller inre vattenvägar ( C5-0208 / 1999 - 1998 / 0106 ( COD ) ) ( föredragande : Koch ) Herr talman , mina damer och herrar !
Beträffande den andra behandlingen kan kommissionen bara godkänna ett ändringsförslag som föreslagits av parlamentet .
Detta förslag tar kommissionen upp och godkänner .
( Talmannen förklarade den gemensamma ståndpunkten godkänd ( efter dessa ändringar ) . )
Betänkande ( A5-0104 / 1999 ) av Koch för utskottet för regionalpolitik , transport och turism om förslaget till Europaparlamentets och rådets direktiv om ändring av direktiv 94 / 55 / EG om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg ( KOM ( 1999 ) 0158 - C5-0004 / 1999 - 1999 / 0083 ( COD ) ) ( Parlamentet antog lagstiftningsresolutionen . )
Betänkande ( A5-0108 / 1999 ) av Schroedter för utskottet för regionalpolitik , transport och turism om meddelandet från kommissionen - Strukturfonderna och samordningen med Sammanhållningsfonden - Riktlinjer för programmen för perioden 2000-2006 ( KOM ( 1999 ) 0344 - C5-0122 / 1999 - 1999 / 2127 ( COS ) ) ( Parlamentet antog resolutionen . )
Betänkande ( A5-0107 / 1999 ) av Berend för utskottet för regionalpolitik , transport och turism om den sjätte periodiska rapporten om den sociala och ekonomiska situationen i Europeiska unionens regioner ( SEK ( 1999 ) 0066 - C5-0120 / 1999 - 1999 / 2123 ( COS ) ) ( Parlamentet antog resolutionen . )
Betänkande ( A5-0069 / 1999 ) av von Wogau för utskottet för ekonomi och valutafrågor om kommissionens vitbok om modernisering av reglerna om tillämpning av artiklarna 85 och 86 i EG-fördraget ( KOM ( 1999 ) 0101 - C5-0105 / 1999 - 1999 / 2108 ( COS ) ) ( Parlamentet antog resolutionen . )
Betänkande ( A5-0078 / 1999 ) av Rapkay för utskottet för ekonomi och valutafrågor om den XXVII : e rapporten om konkurrenspolitiken - 1998 ( SEK ( 1999 ) 0743 - C5-0121 / 1999 - 1999 / 2124 ( COS ) ) ( Parlamentet antog resolutionen . )
Betänkande ( A5-0087 / 1999 ) av Jonckheer för utskottet för ekonomi och valutafrågor om den sjunde översikten över statligt stöd i Europeiska unionen inom tillverkningsindustrin och vissa andra sektorer ( KOM ( 1999 ) 148 - C5-0107 / 1999 - 1999 / 2110 ( COS ) ) ( Parlamentet antog resolutionen . )
Betänkande ( A5-0073 / 1999 ) av Langen för utskottet för ekonomi och valutafrågor om kommissionens rapport om 1998 års genomförande av kommissionens beslut nr 2496 / 96 / EKSG av den 18 december 1996 om gemenskapsregler för statligt stöd till stålindustrin ( gemenskapsreglerna för stöd till stålindustrin ) ( KOM ( 1999 ) 94 - C5-0104 / 1999 - 1999 / 2107 ( COS ) ) ( Parlamentet antog resolutionen . )
Röstförklaringar- Egna medel Europeiska unionen finansieras uppenbarligen med fyra slags egna medel .
Men den europeiska budgeten grundas i själva verket på moms och BNI-uttag , framför allt sedan man övergav gemenskapspreferensen och flerfaldigade antalet frihandelsområden , och därigenom urholkade tullavgifterna och den gemensamma jordbruksskatten , vilka redan har decimerats av de allmänna preferenssystemen .
Bedrägerier i fråga om gemenskapsmomsen och felaktiga beräkningar av BNI , som är det fjärde medlets beskattningsbara bas , påverkar i känsliga proportioner gemenskapens medel , såväl intäkterna som ur rättvisesynpunkt .
Det Europa som när federala anspråk finansieras därmed mer än någonsin som den enkla mellanstatliga organisation det egentligen är , men som det vägrar att vara .
Det framgår tydligt i den förordning vi nu behandlar .
Här ägnar man sig åt " bokföringen av de egna medlen " , " tillhandahållandet " av dem och över " kontrollen " av de fastställda rättsenliga belopp som ställts till kommissionens förfogande .
I den nyinrättade rådgivande kommittén ingår dessutom företrädare från de skattebetalande medlemsstaterna .
Här är det långt till avarter som en " gemensam straffrätt " , en " gemensam allmän åklagare " eller gemenskapspolis , i och med OLAF .
Här finns det ännu ingen europeisk federal skatt .
Men det stämmer att ett Europa med 25 medlemmar fordrar en europeisk inkomstskatt , om det nu inte blir vinster som kommer att beskattas , eller en koldioxidskatt som finansierar 2025 års budget .
Betänkande ( A5-0105 / 1999 ) av Koch Det är med stor tillfredsställelse jag välkomnar detta betänkande om en bättre harmonisering inom utbildningen av säkerhetsrådgivare för transport av farligt gods .
Under de senaste åren har de nationella och internationella transporterna av farligt gods ökat avsevärt , vilket har ökat olycksriskerna .
Vissa av olyckorna har berott på en otillräcklig kunskap om de risker som hänger samman med den här typen av transporter .
Det har således visat sig nödvändigt att anta åtgärder - inom ramen för genomförandet av den inre marknaden - för att ombesörja ett bättre förebyggande av risker .
Genom direktiv 96 / 35 / EG uppfylldes det kravet .
Följaktligen har de företag som transporterar farligt gods och de företag som genomför lastning och lossning i samband med sådana transporter med rätta sett sig tvingade att respektera regler om riskförebyggande , vare sig det gäller transporter på väg , järnväg eller inre vattenvägar .
För att göra det lättare att förverkliga detta mål , föreskrev direktiv 96 / 35 / EG att de säkerhetsrådgivare som utses för transporter av farligt gods skall ha en lämplig yrkesutbildning .
Målet med denna yrkesutbildning för rådgivare skulle vara en kunskap om de viktigaste lagar , förordningar och bestämmelser som gäller för dessa transporter .
Detta utgjorde ett framsteg för några år sedan , men så småningom uppstod problem eftersom det saknas specifika bestämmelser om harmoniseringen av examineringsvillkoren .
Det föreföll därför nödvändigt att komma tillrätta med den svagheten , för att nå en högre och enhetlig utbildningsnivå för säkerhetsrådgivare , men också för att undvika skillnader mellan utbildningskostnader och följaktligen en inverkan på konkurrensen mellan medlemsstaternas företag .
Kommissionens förslag syftar till att garantera en enhetlig utbildning av säkerhetsrådgivarna .
Förslaget avgränsar minimiinnehållet i en examen och fastställer den behöriga myndighetens uppgifter , såväl som vilka krav som skall uppfyllas av examineringsorganen .
Parlamentet har ställt sig positivt till denna text .
Men det har ändå lagt fram flera ändringsförslag , varav de flesta har införlivats i rådets gemensamma ståndpunkt , t.ex. att det skall vara nödvändigt att genomföra en fallstudie och ge utlåtande om tillstånd till vissa dokument inom ramen för en " specificering av de examineringsformer som examineringsorganet föreslår " .
Jag ger för övrigt mitt stöd till att tidsfristen för genomförandet av dessa bestämmelser skjuts upp till tre månader efter det att direktivet har trätt i kraft , med hänsyn till vad som är realistiskt .
Jag vill avsluta genom att insistera på det faktum att rådgivarnas yrkeskvalifikationer kommer att bidra till en förbättrad servicekvalitet till användarnas fördel , och det kommer att minimera de olycksrisker som en försämrad miljö kan medföra liksom de allvarliga skador vilka kan skada den fysiska integriteten hos alla de personer som kan komma i kontakt med farligt gods .
Betänkande ( A5-0104 / 1999 ) av Koch I oktober förra året uttalade jag mig om Hatzidakisbetänkandet om transport av farligt gods på järnväg .
Mina synpunkter i dag står inte långt ifrån dem jag hade då .
De kan sammanfattas på följande sätt : jag beklagar att vi ständigt skjuter upp antagandet av harmoniserade normer på ett så avgörande område som transport av farligt gods .
Det skadar människors säkerhet och miljön .
Jag vill erinra om att ett direktiv om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg trädde i kraft den 1 januari 1997 .
Det innehåller ett antal övergångsbestämmelser som var giltiga fram till den 1 januari 1999 .
Från och med det datumet borde vi ha uttalat oss om ett förslag från Europeiska kommissionen , med syftet att få dessa undantag att upphöra .
Enligt det nuvarande förfarandet är det Europeiska standardiseringskommittén ( CEN ) som föreslår normer på det här området .
Dessa upptas sedan i Europeiska överenskommelsen om internationell transport av farligt gods på väg , som undertecknades i Genève 1957 ( mer känt under förkortningen ADR ) och tillämpas i hela Europa , och vars bestämmelser utgör grunden för den lagstiftning som är tillämplig i Europeiska unionen .
Men CEN har inte kunnat utföra sitt arbete inom den anvisade tiden .
Syftet med det förslag från kommissionen som vi diskuterar i dag är därför att ändra på direktivet för att lösa problemen på kort sikt , och inte att sätta punkt för övergångssystemet , vilket borde ha varit fallet !
Precis samma sak hände när det gällde transport av farligt gods på järnväg , fast med en skillnad : en tidsfrist fastställdes .
I dag har vi inte den blekaste aning om när CEN kommer att kunna ge oss konkreta förslag .
Fram till dess är det egentligen onödigt för medlemsstaterna att ändra sina nationella bestämmelser .
I betänkandet accepteras också att man inför en viss flexibilitet , och man tillerkänner staterna möjligheten att anta eller tillämpa olika normer .
Medlemsstaterna skulle således kunna fortsätta att tillämpa sina egna normer för vissa transportabla tryckbärande anordningar , eftersom de europeiska normerna inte är tillräckliga i det fallet .
Staterna kan också anta olika bestämmelser för transporter av lokal art och enstaka transporter .
Med denna röstförklaring vill jag i dag uttrycka mitt djupa missnöje och min stora oro .
Betänkande ( A5-0108 / 1999 ) av Schroedter Herr talman !
Jag skulle vilja lägga tyngd bakom min röstförklaring genom denna muntliga förklaring med anledning av Schroedterbetänkandet om den regionala utvecklingen .
Jag vill uppmana såväl medlemsstaterna som kommissionen att ägna tillräcklig uppmärksamhet åt de stora välfärdsskillnader som finns kvar mellan de olika regionerna i Europa .
Det gäller inte bara skillnaden i inkomst per capita , utan det är framför allt de stora skillnaderna beträffande sysselsättning som fortsätter att vara en källa till oro .
Trots det faktum att gemenskapen , bland annat via strukturfonderna , lägger ned avsevärda summor på att bekämpa skillnaderna mellan chanserna till utveckling för våra regioner i Europa kvarstår dessa skillnader .
Det gör att jag ställer mig frågan om inte gemenskapen bör lägga om kursen på ett mer drastiskt sätt , och på grundval av mycket strikta utvärderingar bör övergå till en kursändring och till en ändring av målsättningarna som gör det möjligt att bedriva en effektivare kamp mot skillnaderna i välfärd och sysselsättning .
Herr talman !
Vad gäller Schroedters betänkande är jag medveten om , och har fått bekräftat av Barnier , att reglerna om komplementaritet vad strukturfonderna beträffar bara kan tillämpas på medlemsstatsnivå och inte är tillämpliga på ett transitivt och öppet sätt inom medlemsstaterna till förmån för självstyrande regioner såsom Wales eller Skottland .
Jag tycker att detta är mycket otillfredsställande .
Jag hoppas att vi kan ompröva denna fråga vid ett senare tillfälle .
Jag vill göra klart att jag har denna viktiga invändning även om jag röstade för betänkandet . .
( EN ) I Schroedters betänkande talar man om behovet att främja partnerskap vad beträffar ianspråktagandet av EU : s strukturfonder för perioden 2000-2006 .
Jag anser att detta är särskilt viktigt eftersom medlen i EU : s strukturfonder alltid används på ett sätt som maximerar olika regioners ekonomiska utveckling när lokala och regionala myndigheter är involverade i beslutsfattandet om hur dessa fonder skall användas .
I egenskap av ledamot av Europaparlamentet för Leinsters valkrets har jag alltid hävdat behovet av att förverkliga lokala initiativ som stöds av nationella EU-fonder .
Jag anser att den irländska regeringen och Europeiska kommissionen och olika EU-regeringar inte själva kan besluta om specifika utgiftsprioriteringar .
Jag anser att lokala myndigheter och grupper från den privata sektorn och frivilligsektorn bör vara fullt involverade i beslutsfattandet om hur de europeiska strukturfonderna skall användas .
Vi har till exempel sett vilken framgång programmen Leader I och II har haft i Irland i form av de arbeten som har skapats genom dessa program på den irländska landsbygden och inom Europa .
Programmet Leader III skall verkställas någon gång senare i år .
Kärnan i Leader-programmet är att ge offentliga , privata och ideella grupper möjlighet att slå ihop sina resurser så att en permanent och hållbar sysselsättning skapas i små och medelstora företag på landsbygden .
Detta är ett klassiskt exempel på hur partnerskapskonceptet fungerar , och sådana program måste ingå i dess befogenheter .
Den europeiska fonden för fred och försoning har också varit framgångsrik när det gäller att skapa arbetstillfällen i Irlands gränsområden .
Även här finns ett aktivt deltagande från offentliga , privata och ideella grupper vilka lämnar förslag om hur särskilda fondmedel bäst kan användas för att understödja olika lokala projekt för att skapa sysselsättning i denna region .
Under nästa runda för EU : s strukturfonder 2000-2006 kommer andra EU-initiativ såsom " Equal " och " Urban " att vara i full gång .
Dessa initiativ måste också involvera för att identifiera var de europeiska strukturfonderna kommer bäst till nytta .
Föredraganden hänvisar till behovet att skapa en samordnad inställning till planer och program för nya EU-strukturfonder .
De måste främja ett decentraliserat , effektivt och mångsidigt partnerskap grundat på kunskaperna och engagemanget inom regionala och lokala myndigheters alla sektorer .
Detta är mycket känsligt eftersom avgörande ekonomiska och sociala problem i vårt land inte kan lösas om det inte finns en samordning av nationell , europeisk och lokal bidragsgivning .
Detta betänkande föranleder följande fråga : vilket är regionalpolitikens existensberättigande ?
För att minska de regionala skillnaderna givetvis .
Men det hänger framför allt samman med den europeiska marknaden , som a priori skall garantera oss en bättre fungerande ekonomi , men som också kan vara en källa till orättvisor .
Jacques Delors brukade säga att marknaden är närsynt , därav den politiska nödvändigheten av att minska skillnader .
Det handlar om den solidaritet som är ursprunget till den europeiska sociala modell som vi alla försvarar , och som har gett upphov till den ekonomiska och sociala sammanhållningen .
Det verkliga politiska målet , på samma sätt som när det gäller ekonomi och valutafrågor , är något som utvecklas i samarbete med medlemsstaterna , regionerna och de lokala myndigheterna .
Kommissionens uppgift är att med hjälp av riktlinjer visa medlemsstaterna vilken linje som skall följas , för att de eftersträvade målen skall uppnås inom ramen för programplaneringen .
Därför kommer jag att stödja detta betänkande , samtidigt som jag beklagar , av skäl som har att göra med tidsplanen , att Europaparlamentet inte rådfrågades förrän mycket sent i fråga om de riktlinjer som skall hjälpa medlemsstaterna , regionerna och de lokala myndigheterna med programplaneringen av mål 1 , 2 och 3 .
I övrigt önskar jag att kammaren också tar hänsyn till yttrandet från utskottet för sysselsättning och sociala frågor , vilket tillfogar en reflektionsplan för centrala frågor såsom bekämpningen av social utslagning , stödet till den sociala ekonomin och genomförandet av sysselsättningsstrategin .
Schroedters arbete är ett steg mot en större öppenhet och effektivitet inom ramen för de strukturella stöden .
Hon sätter värde på den växande och ytterst viktiga roll som samtliga aktörer har , och särskilt våra lokala partner - de enda som kan definiera specifika frågor och sociala problem .
Därför vill vi försäkra oss om att de partnerskap som skall genomföras blir verkliga partnerskap , decentraliserade partnerskap som involverar samtliga berörda aktörer , och därför omformulerar vi vårt krav på att det skall inrättas ett centrum för förvaltning av strukturstöden i medlemsstaterna , med uppdraget att samordna genomförandet och förvaltningen av stöden .
För det ändamålet krävs det att utvärderingskommittéerna står öppna för Europaparlamentets ledamöter , föreningar , näringsidkare som berörs av projekten samt det civila samhället .
Dessa riktlinjer är ett steg för att göra gemenskapens strukturstöd effektivare .
Ändras de enligt Schroedterbetänkandet , går de i rätt riktning .
De uppmanar också till en allmän debatt om sammanhållningspolitikens framtid efter år 2006 , men det är en annan debatt .
Låt oss stödja detta första steg i väntan på den . .
( EN ) I detta betänkande krävs drastiska nedskärningar av det illegala statliga stöd vissa medlemsstater delar ut .
Även om jag helhjärtat stöder detta syfte skulle jag mycket hellre se att ett sådant stöd avskaffades helt .
Enligt min mening är illegalt statligt stöd inte mycket bättre än statligt sponsrad social dumpning .
Vi är alla emot social dumpning när förövaren är den välmående bilindustrin , då måste vi också vara emot den när förövaren är en regering .
Om vi skall kunna få en effektiv inre marknad som gör den europeiska industrin konkurrenskraftig globalt och skapar välstånd och sysselsättning för alla européer måste vi ha en jämn spelplan .
Illegalt statligt stöd däremot förstör konkurrenskraftiga företag och skapar arbetslöshet .
Det finns förstås fall där statligt stöd kan vara nödvändigt och legitimt , för att till exempel hjälpa företag vid omstruktureringar .
I alla sådana fall måste dock strikta kriterier uppfyllas och tillstånd från Europeiska kommissionen inhämtas i förväg .
Oavsett om vi talar om nötkött till Frankrike eller mutor till industrin får inte EU : s medlemsstater tillåtas att driva gäck med lagen .
Jag stöder med entusiasm förslaget i betänkandet att offentliggöra en " resultattavla " som visar det statliga stödet per medlemsstat .
Länder som hävdar att de ligger i Europas hjärta men som systematiskt bryter mot dess regler bör demaskeras och deras hyckleri avslöjas .
Medlemsstaterna kan inte tillåtas proklamera europeisk solidaritet offentligt och samtidigt försöka underminera den inre marknaden privat .
Jag blir något uppmuntrad av det faktum att nivån på det statliga stödet till industrin i Europa tycks minska .
Emellertid återstår mycket att göra , och jag uppmanar kommissionen att vara mycket tuffare när den exponerar Europas bidragsnarkomaner . - ( PT ) Eftersom kommissionens viktigaste instrument för att övervinna de regionala skillnaderna är strukturfonderna och Sammanhållningsfonden , är det väsentligt att Europaparlamentet deltar i utformandet av dess allmänna vägledande riktlinjer utan att det sker på bekostnad av subsidiariteten , då fastställande av utvecklingsstrategierna i varje land är medlemsstaternas sak .
Tyvärr har Europeiska kommissionen redan gått framåt med sina riktlinjer och parlamentets ståndpunkt är inte mycket värd för programmen under perioden 2000-2006 .
Det är dock viktigt att trycka på betydelsen av att dessa fonder först och främst prioriterar utvecklingen i de länder och regioner som har störst svårigheter och i gemenskapens yttersta randområden , vilket Portugal och regionerna Azorerna och Madeira är exempel på , för att uppnå ekonomisk och social sammanhållning .
I själva verket uppfyller inte kommissionens riktlinjer dessa mål helt .
Det är också viktigt att det finns precisa indikationer och tillräckliga medel för att skapa kvalitativ sysselsättning med rättigheter liksom för att effektivt främja lika rättigheter och möjligheter , stödja en social och solidarisk ekonomi , landsbygdens utveckling , de små och medelstora företagarna , samt för att förbättra livskvaliteten för stadsbefolkningen i fattigare områden , främst inom området för bostäder som subventioneras med allmänna medel , för att härigenom uppnå en hållbar utveckling i städerna . .
( IT ) Om innehållet i artikel 158 i EG-fördraget syftar till att främja en harmonisk utveckling av hela gemenskapen , så måste vi tyvärr konstatera att vi fortfarande är långt från målet att utjämna skillnaderna .
Det är till och med så , till exempel för de italienska områden som återförts till mål 1 , att skillnaderna paradoxalt nog ökar , framför allt på grund av att de lokala organisationernas förmåga att hantera gemenskapens rutiner fortfarande är bristfällig och att det råder ett permanent kaos när det gäller förvaltningen .
Trots ingreppen i regelsystemet har vi ännu inte lyckats få gemenskapens strukturer att arbeta snabbare .
Om man inte förenklar byråkratin så blir det svårt att uppnå gemenskapens mål , som är att genomföra reformer präglade av effektivitet och koncentration .
I det avseendet är kommissionens dokument bristfälligt , eftersom här inte finns några som helst rekommendationer till medlemsstaterna om hur man skall kunna förenkla nationella regler och rutiner när det gäller hur de nationella myndigheterna skall presentera och informera om olika projekt , eller när det gäller finansiering , genomförande och kontroll .
Små och medelstora företag , mikroföretag och hantverkare är fortfarande " svaga subjekt " , eftersom de hinder som finns i regler och byråkratiska rutiner i vissa medlemsstater , bland annat Italien , just för dem gör det betydligt svårare att få tillgång till strukturfonderna .
Ett viktigt handicap är regionernas och andras oförmågan och bristande möjligheter att planera i god tid , varför kommissionen , som på grundval av beslutet om riktlinjer 97 / 99 ( Howittsbetänkandet ) hade kunnat rådfråga parlamentet i god tid , i själva verket hittade ett bekvämt alibi när man inrättade den förkortade planeringsfasen i medlemsstaterna och offentliggjorde riktlinjerna redan i juli 1999 , dvs. innan det nyvalda parlamentet hade inlett sitt arbete .
På det viset hindrade man parlamentet att påverka riktlinjernas utformning .
Av den anledningen blir halvtidsbedömningen av artikel 42 i förordningen 1260 / 99 betydelsefull .
De nuvarande riktlinjerna utmärks generellt sett inte av klarhet och öppenhet .
Trots att det är en viktig fråga berör de bara ytligt möjligheten att mäta de framsteg som gjorts utifrån verifierbara mål och i enlighet med gemenskapspolitikens strategier , och man uppehåller sig inte i tillräckligt hög grad vid utvidgningens effekter , och inte heller innehåller riktlinjerna specifika föreskrifter eller förtydliganden i frågan , vare sig för de regionala och nationella myndigheterna eller för kandidatländerna .
Men oavsett detta är vi trots allt positiva till att man i riktlinjerna ställer de geografiska målen åt sidan och riktar in sig på sektoriell politik .
Även om detta , teoretiskt sett , kan uppfylla kravet på koncentration och därmed kravet att åtgärderna skall vara effektiva , så uppkommer spontant frågan om den nuvarande situationen i mål 1-området är sådan att den faktiskt gör en integrerad politik möjlig .
För att fullfölja en sådan skulle det krävas ett operativt samordnande instrument för avsättningarna .
Vi kan därför , i princip , ge ett positivt svar på kommissionens begäran att få inrätta ett centrum för att främja strukturen i medlemsstaterna , men enbart genom att samordna förverkligandet och genomförandet av strukturella insatser på plats , så att ett sådant centrum inte blir till ett instrument för centralisering på övernationell nivå och att det garanterar att uppmärksamheten verkligen riktas mot de områden - jag säger det ännu en gång - som på grund av ett antal samverkande negativa faktorer ännu inte har nått upp till rätt nivå när det gäller att utnyttja strukturfonderna , för annars skulle det faktum att man ersätter det geografiska målet med sektorpolitik kunna sluta i en åtgärd som i själva verket blir negativ .
Riktlinjerna innebär , i det skick de godkänts av kommissionen , en allvarlig begränsning eftersom de i stället för att uppfylla syftet att ange en inriktning räknar upp en katalog av tänkbara föreskrifter , en katalog som , eftersom den inte är prioriterad , i själva verket skulle kunna få medlemsstaterna att gå vilse genom att rikta deras uppmärksamhet mot ett brett urval av olika förslag , vilket skulle stå i strid mot den önskvärda koncentrationen .
Vi skulle kunna säga att det verkar som om man ännu en gång har förlorat en chans att effektivt verka för en hållbar utveckling i städerna genom att bromsa den tilltagande urbaniseringen och den därmed följande förstöringen av landskapet .
Man har inte i tillräckligt hög grad tagit hänsyn till betydelsen av generella subventioner , något som skulle kunna visa sig mycket användbart för att återskapa en balans mellan stad och land och dessutom vill man inte ge de lokala myndigheterna rätten att självständigt bestämma villkoren för en utveckling av sina territorier på kort sikt och genom egna åtgärder bidra till strukturfondernas reformansträngningar och till att målen effektivitet , koncentration och en snabbare byråkrati uppnås .
Landsbygden måste äntligen betraktas som en tillgång som vi hela tiden måste investera mera i så att vi ger ungdomarna en anledning att stanna på landsbygden för att på så vis undvika att den faller sönder ekonomiskt och socialt .
Det är ett numera välkänt faktum att för att uppnå det målet måste man i landsbygdsområdena skapa arbetstillfällen som inte bara är knutna till det traditionella jordbruket - även om det också är viktigt för att skydda miljön och den biologiska mångfalden - utan snarare inom sektorer som turism , idrott , kultur , miljö , små och medelstora företag , tjänster .
Ett verkligt tomrum finns det i riktlinjerna på grund av bristen på konkreta förslag för att förverkliga samordningen mellan strukturfonderna och en strategi för ökad sysselsättning , en samordning som , just därför att den tillämpas för första gången under programperioden 2000-2006 , förutsätter att medlemsstaterna har behov av " riktlinjer " .
Det bör även understrykas att kommissionen ännu en gång undviker problemet med konkreta åtgärder inom området lika möjligheter .
Slutsatsen blir att detta är ett dokument som inte är särskilt tillfredsställande och i vissa avseenden en ren besvikelse .
Betänkande ( A5-0107 / 1999 ) av Berend - ( PT ) Vi stöder i det väsentliga den bedömning och de överväganden föredraganden gör angående den sjätte periodiska rapporten om den sociala och ekonomiska situationen och utvecklingen i Europeiska unionens regioner .
Vi begränsar oss därför till att betona några aspekter .
För det första , och som kommissionen själv säger , berodde de kraftiga framstegen i BNI per capita i vissa fattiga regioner mellan 1991 och 1996 i hög grad på att de nya tyska delstaterna togs med i beräkningarna av gemenskapens genomsnitt , från första året , vilket var uppenbart avgörande för den påtagliga minskningen av unionens BNI per capita .
Därefter anser vi det vara av särskild betydelse att konstatera att återhämtningen som har skett i vissa regioner åtföljdes av en mycket liten ökning av sysselsättningen , något som därför kräver nya utvecklingsstrategier , med ett mycket större engagemang inom detta område .
Denna situation talar emot en minskning av sysselsättningsskapande åtgärder till enbart medlemsstaterna , såsom föreslås i rapporten .
Sist men inte minst , en hänvisning till föredragandens förslag om att denna typ av rapporter i framtiden , bland andra aspekter , också skall innehålla en analys av hur sammanhållningen mellan regioner i varje land utvecklas .
Den mängd olika situationer och olika utvecklingsmönster som region för region uppvisas inom samma land , kräver i själva verket en fördjupad analys av denna fråga som gör det möjligt att förändra regionalpolitiken ( eller andra politikområden ) för att garantera sammanhållningen också inom varje medlemsstat .
Berendbetänkandet erbjuder oss en intressant analys av den ekonomiska situationen och utvecklingen i Europeiska unionens regioner .
Men den franska delegationen i Gruppen Unionen för nationernas Europa tar avstånd från vissa av de påståenden som finns i betänkandet .
Punkt 26 " påpekar att det särskilt behövs en konsolidering av budgeten såsom förutsättning för att den ekonomiska och monetära unionen och utvidgningen av unionen skall kunna genomföras med framgång " .
När medlemsstaterna är förpliktade att genomgå en strikt finansiell bantningskur för att uppfylla konvergenskriterierna - det var för övrigt berättigat att de själva ansträngde sig för det - ger federalisterna prov på en mycket förvånande ekonomisk glupskhet .
För att visa att man erkänner EMU : s och sammanhållningspolitikens misslyckande , säger man att bristen på uppnådda resultat beror på en brist på pengar .
Alla tävlar vältaligt om att kräva mer medel , men det finns ingen som funderar på om de utbetalade pengarna är effektiva .
Vad skall man säga om ett budgetförfarande som går ut på att fastställa utgiftsmål i stället för utgiftstak , att - kosta vad det kosta vill - söka efter projekt för att med alla krafter spendera de anslagna medlen , i stället för att bevilja medel till befintliga projekt ?
Utgiften blir ett mål i sig och ett bevis på att ett program har lyckats .
Den statistik som Europeiska kommissionen offentliggör i sin sjätte översikt visar trots allt , vilket Berend underströk , den förda politikens begränsningar .
Europeiska unionens rikaste regioner har ökat i betydelse mellan 1986 och 1996 , vilket vittnar om att rikedomar , arbetstillfällen och aktiviteter har koncentrerats till vissa områden : Hamburg , Bryssel , Anvers , Luxemburg , Ile-de-France , Darmstadt , Oberbayern , Bremen , Wien , Karlsruhe och Emilia-Romagna .
I motsats till vad föredraganden hävdar , kommer Ekonomiska och monetära unionen att bidra till flykten från de mest avlägsna , mest lantliga och minst befolkade regionerna , till förmån för unionens centrala linje ( Benelux , nordvästra Tyskland , Norditalien , Île-de-France ... ) .
De fattigaste regionerna kommer steg för steg i kapp utvecklingsmässigt .
Genomsnittet för de tio fattigaste regionerna uppnådde 41 procent av gemenskapens BNP år 1986 .
År 1996 låg det på 50 procent .
Framstegen är särskilt tydliga i Portugal och Irland .
Om de rikare blir allt rikare och de mycket fattiga blir mindre fattiga , verkar det som om genomsnittsregionerna , de som lyder under mål 2 , i realiteten har fått en lägre BNP , i vissa fall en icke försumbar minskning , samt försämrade sysselsättningsförhållanden .
Det är särskilt tydligt i Frankrike : i regionen Champagne-Ardennes , som jag har den äran att företräda , har BNP minskat från 105 till 94 procent av EU-genomsnittet , i Pays-de-Loire har den sjunkit från 95 till 91 procent , i Auvergne från 89 till 83 procent .
Detta är en generell tendens , som varken besparar Rhône-Alpes eller Alsace .
Den bekräftas i Sverige och Finland , länder där arbetslösheten under de senaste åren har ökat i oroande proportioner , liksom i flera av Förenade kungarikets regioner .
Därför kan det tyckas märkligt att mål 2 - vilket anslås till industri- och landsbygdsregioner som genomgår en ekonomisk omstrukturering - offrades i reformen av strukturfonderna till förmån för mål 1 och 3 : för perioden 1999-2006 ligger dess totalanslag på 22,5 miljarder ecu , en siffra som i princip är densamma som för perioden 1994-1999 .
De landsbygdsregioner som är berättigade till mål 5b kan räknas till de främsta offren för denna situation : i Frankrike kommer 27 procent av den befolkning som är berättigade till strukturfonder att förlora sin rätt vid övergångsperiodens slut .
Denna siffra är mycket högre i vissa regioner , såsom Pays de la Loire , Alsace och Basse-Normandie , högerns väljarbastioner som fallit offer för den pluralistiska vänsterregeringens politiskt förslagna klientilism .
Med stöd av sådana beslut är det tveksamt om regionalpolitiken kan bidra till en harmonisk fysisk planering i Europeiska unionens medlemsstater .
Betänkande ( A5-0069 / 1999 ) av von Wogau Med hänsyn till sysselsättningsläget i gemenskapen och Europeiska unionens uttalade ambition att resolut bekämpa arbetslösheten , bör kommissionens analys av koncentrationer ta hänsyn till andra faktorer än konkurrensen .
Som ett exempel skall jag ta upp företaget ABB-Alsthom Power , som har en stor delegation anställda från hela Europa närvarande i dag i Strasbourg .
Ledningen i ABB-Alsthom Power , ett resultat av en fusion som genomfördes i juni 1999 , har tillkännagivit en omstrukturering som redan nu innebär att arbetstillfällen kommer att avvecklas i ett antal länder .
Denna ödesdigra situation för sysselsättningen föranleder flera frågor , bl.a. om vilken information som har tillhandahållits det europeiska företagsrådet , som har funnits sedan 1996 .
Och det förutsätter en förnyelse och förstärkning av gemenskapens direktiv om europeiska företagsråd .
Det förutsätter också en kontroll av koncentrationer , vilken skall ta hänsyn till sysselsättningen , miljön och konsumenterna .
Eftersom betänkandet från utskottet för ekonomi och valutafrågor är otillräckligt ur den synvinkeln , har jag avstått från att rösta . - ( PT ) När kommissionen försöker tillämpa subsidiaritetsprincipen på gemenskapens konkurrenspolitik , decentraliserar man ansvaret för beslut och missbruk av dominerande ställning vad gäller företagsavtal som skapar snedvridning på marknaden , till nationella myndigheter och domstolar även om de fortfarande hör till anmälningssystemet för frågor om företagskoncentration och statligt stöd .
Den ståndpunkt som nu har intagits är en strävan att skapa snabbare och billigare former för tillämpningen av konkurrenspolitiken , genom att EG-rätten tillämpas av de nationella domstolarna och inte av EG-domstolen , och även en inriktning mot specialdomstolar .
Denna partiella åternationalisering av konkurrenspolitiken kan medföra ökade kostnader för medlemsstaterna .
Å andra sidan , vilket föredraganden erinrar om , har ofta statliga monopol , i konkurrenspolitikens namn bytts ut mot privata monopol med privatisering av viktiga statliga sektorer och företag , så som är fallet i Portugal , med negativa följder för landet och för dess arbetare .
Kommissionens vitbok om en modernisering av reglerna om tillämpning av artiklarna 85 och 86 i EG-fördraget ( de nya 81 och 82 ) föreslår självklart inte en " åternationalisering " av konkurrenspolitiken , vilket vissa i Europaparlamentet fruktar .
Men den låter ana ganska intressanta utvecklingsmöjligheter för Europeiska unionen .
Kommissionen konstaterar att dess enheter översvämmas av förhandsanmälningar om avtal mellan företag som skulle kunna snedvrida konkurrensen , och fruktar att de kommer att bli fler när nya medlemmar tillkommer .
Den föreslår därför att man avskaffar det nuvarande systemet , dvs. att dessa avtal skall godkännas i förväg , och att tillämpningen av konkurrensreglerna skall decentraliseras till medlemsstatsnivå .
Det mest anmärkningsvärda är enligt min mening den signal som detta förslag ger oss : kommissionen föregriper utvidgningens konsekvenser och anser att den med nödvändighet , ja nästan med automatik , förutsätter en reform av det centraliserade systemet .
Denna reform består givetvis i en uppmjukning och inte en nedmontering .
På papperet skall kommissionen behålla kontrollen och den centrala ledningen i det nya systemet .
Betänkandet av von Wogau , som Europaparlamentet just har röstat igenom , uppmuntrar för övrigt kommissionen på den punkten .
Men samtidigt kan man lätt se att det sammanbrott som utvidgningen medför kan leda till en begränsning av gemenskapens behörigheter , och till en utvidgad subsidiaritet .
Det är ett annat Europa som på sikt kan komma att ta form .
Är det förresten inte just det som skrämmer vissa socialister i Europaparlamentet ?
De tyska socialdemokraterna röstade emot betänkandet av von Wogau , eftersom de anser att det skulle sönderdela den europeiska konkurrenspolitiken , i klartext skada den likriktande överstaten .
Märkligt nog har ett arbetsgivarparti anslutit sig till dem , eftersom det föredrar det europeiska systemet med " en enda lucka " , vilket för dem verkar vara mer ekonomiskt och mer stabilt juridiskt sett .
Det är faktiskt en fördel med det nuvarande systemet .
Men ur en annan synvinkel bör man också betänka att starten av den decentralisering som inleds i dag på sikt kan leda till en större frihet när det gäller hänsynstagandet till varje lands behov , något som kommer alla till del .
Betänkande ( A5-0078 / 1999 ) av Rapkay De förtroendevalda i Lutte Ouvrière kommer inte att rösta för dessa betänkanden om den europeiska konkurrenspolitiken .
Konkurrensen , dvs. det krig som de stora företagen för sinsemellan , tar sig ständigt uttryck i uppsägningar , nedläggningar av företag , för att inte tala om ett oändligt slöseri när det gäller utnyttjandet av den produktiva kapaciteten .
Vi har fått ytterligare ett exempel på detta i och med att trusten ABB Alsthom Power kommer att avveckla arbetstillfällen i Europa .
18 miljoner arbetslösa , 50 miljoner fattiga i Europeiska unionen , som trots allt är en av de rikaste regionerna i världen : däri ser vi resultatet av den konkurrens som EU-institutionerna har för avsikt att främja .
Kommissionens vilja att reglera konkurrensvillkoren på den europeiska marknaden är löjeväckande , för den enda lag som konkurrensen lyder under är djungelns lag , dvs. att de mäktigaste krossar eller slukar de svagaste .
Det är upprörande , framför allt ur en social synvinkel .
Europeiska kommissionens rapport visar utan omsvep att unionens institutioner endast intresserar sig för de stora kapitalistiska företagsgrupperna , som hänger sig åt detta ekonomiska krig och inte på något sätt åt de offer som de själva skapar .
Ingenting för att förhindra arbetslöshetens utbredning , ingenting för att skydda löntagarna , ingenting för att förhindra att de stora företagen driver en del av befolkningen till armod enbart för att skapa ännu större rikedomar för sina aktieägare !
Skall vi medge att det finns en fördel med denna rapport , är det att den visar för samhällets arbetande majoritet att den inte kan hoppas på att EU-institutionerna kommer att upprätthålla , och än mindre förbättra deras levnadsvillkor . - ( PT ) När föredraganden uttalar sig om kommissionens årliga rapport om konkurrenspolitiken , påminner han om att konkurrenspolitiken inte kan separeras från social- och miljöpolitiken , utan bör bidra till full sysselsättning , ekonomisk och social sammanhållning , miljöskydd och konsumentskydd .
När föredraganden diskuterar vissa väsentliga instrument för att uppnå de nämnda målen begränsar han sig emellertid praktiskt taget till att kritisera vissa aspekter av de otillåtna statliga stöden och att kräva en harmonisering av bestämmelserna om återbetalning av otillåtna statliga stöd , och ifrågasätter därigenom rätten för de ekonomiskt och strukturellt svagaste medlemsstaterna att stödja ekonomiska sektorer som blivit offer för avreglering och internationell konkurrens .
Å andra sidan ignorerar föredraganden de främsta orsakerna till snedvridningen av konkurrensbestämmelserna , nämligen : den ökade företagskoncentrationen och dess konsekvenser för snedvridning av konkurrensbestämmelserna ; förvandlingen av statliga företag till privata monopol med allvarliga sociala följder , framför allt för sysselsättningen och priset för offentlig service ; olika monopolistiska gruppers missbruk av dominerande ställning genom oacceptabla metoder på miljöområdet och det sociala området , inklusive uppsägningar av tusentals arbetare .
Därav vår röst emot detta betänkande .
Genom att rösta emot detta betänkande gör vi oss till talesmän för alla dem som , i Seattle och överallt i Europa , har markerat sitt motstånd till en värld som reduceras till en strikt handelslogik .
Vi röstar mot detta betänkande med omsorg om utvecklingen av de allmännyttiga tjänsterna , och i synnerhet till minne av offren för tågolyckan i Paddington .
Deras död var inte ett olycksöde utan berodde på en absurd iver att konkurrensutsätta det som borde regleras .
Detta betänkande är i grunden en lågt stående text , som endast inspireras av djungelns lag , för konkurrens kan inte lösa något av de problem som mänskligheten står inför vid detta sekelskifte .
Vare sig det handlar om balansen i biosfären , att främja kulturen eller samarbeta med tredje världen , är en överdriven konkurrens en faktor som hänger samman med tillbakagång och osäkerhet .
Och de 18 miljoner arbetslösa i Europa , tror ni att de är offer för en alltför blygsam tillämpning av konkurrenspolitiken ?
Vi är övertygade om motsatsen , och vi anser inte heller att de statliga stöden per definition är för stora .
Enligt vilken dogm eller vilka effektivitetskriterier skulle de vara för stora ?
Anser ni slutligen att det efter Seattle är seriöst att förespråka en utvidgad roll för WTO ?
Endast de multinationella bolagens juridiska rådgivare kan ge prov på en sådan envishet .
Betänkande ( A5-0087 / 1999 ) av Jonckheer Jag gläder mig åt kvaliteten på den sjunde översikten över statliga stöd i EU och att den numera publiceras årligen , samt åt det faktum att generaldirektoratet för konkurrens använder sin webbplats för att ge både övergripande och mer detaljerad information till allmänheten .
Jag tycker att föredraganden har en bra syn på statliga stöd , och jag vill gratulera honom till det .
Man tenderar alltför ofta att sammanblanda statliga stöd med åtgärder som snedvrider konkurrensen .
Visserligen är en effektiv konkurrenspolitik en förutsättning för att den inre marknaden och den ekonomiska och monetära unionen skall fungera väl .
Samtidigt är den här typen av stöd ibland nödvändiga , vilket föredraganden betonar , och bidrar inte bara till att särskilda företag kan överleva , utan också till en hållbar utveckling ( artikel 6 i fördraget ) , tjänster av allmänt intresse ( artikel 16 ) samt ekonomisk och social sammanhållning ( artikel 158 ) .
Det är likväl uppenbart att stöden måste kontrolleras , ett uppdrag som åligger Europeiska kommissionen .
De stöd som unionens medlemsstater varje år anslår till de granskade sektorerna uppgick till totalt 95 miljarder euro under perioden 1995-1997 , varav 40 procent till tillverkningssektorn .
Det är en avsevärd minskning i förhållande till den föregående perioden , 1993-1995 ( en minskning på 13 procent av det totala beloppet och en minskning från 3,8 till 2,6 procent av stöden till tillverkningssektorn ) .
De minskade stöden kan huvudsakligen förklaras med att stöden till Tysklands nya " länder " har gått tillbaka .
I likhet med föredraganden beklagar jag att de siffror som presenteras i översikten inte täcker samtliga former av statliga stöd .
Europeiska kommissionen bör snarast komma tillrätta med dessa brister .
Den bör också samarbeta med medlemsstaterna för att i god tid förbättra kvaliteten på uppgifterna , dvs. inför den nionde översikten .
Det vore bra om kommissionen offentliggjorde ett register som omfattar beloppen för statliga stöd per medlemsstat .
Jag beklagar också att Europaparlamentet är helt utestängt från den rådgivande kommittén om statliga stöd .
För att kompensera detta bör Europeiska kommissionen lägga fram regelbundna rapporter för oss .
Jag skall avsluta om en aspekt av utnyttjande av statliga stöd som jag tycker verkar särskilt farlig : det gäller de stöd som leder till omlokaliseringar av företag från en medlemsstat till en annan , vilket riskerar att skapa en jakt på subventioner som inte tillför EU : s gemensamma mål någonting .
Därför skulle jag önska att nästa rapport om statliga stöd innehåller en utvärdering av statsstödens effekter på sysselsättningen och mottagarländernas industri och hantverk .
Betänkande ( A5-0073 / 1999 ) av Langen I den viktiga konkurrensdebatten uttalade jag mig i förmiddags om Langens text , som gäller tillämpningen av den sjätte regeln för stöd till stålsektorn under 1998 .
Precis som EG-domstolen slog fast i beslut av den 3 maj 1996 är stålsektorn särskilt känslig för konkurrensrelaterade störningar .
Därför var det berättigat att inrätta ett stödsystem för denna sektor , med ändamålet att garantera de livsdugliga företagens överlevnad , trots att artikel 4 c i EKSG-fördraget förbjuder alla former av statliga stöd till stålsektorn .
Detta är själva syftet med den sjätte regeln om stöd till stålindustrin .
Samtidigt är det givetvis viktigt att förhindra att konkurrensvillkoren kränks och att marknaderna utsätts för allvarliga störningar , varför den här typen av stöd måste regleras .
Det är således nödvändigt att även i fortsättningen begränsa de statliga stöden till att avse forskning , utveckling , miljöskydd samt stöd i händelse av företagsnedläggningar .
På samma sätt är det ytterst viktigt att medlemsstaterna uppfyller sin förpliktelse att till kommissionen anmäla vilka stöd som beviljats deras stålföretag , vilket artikel 7 i de aktuella reglerna föreskriver .
Kommissionen föreslår att staterna skall sända in rapporterna inom två månader efter varje halvårsskifte , och under alla omständigheter en gång per år , utan att kommissionen skall behöva påminna dem om detta .
I likhet med föredraganden gladde jag mig åt kommissionens rapport , men jag beklagade att den inte täcker alla aspekter av statliga stöd .
Även om reglerna för stöd till stålsektorn formuleras på ett mycket tydligt sätt , har kommissionen vid ett flertal tillfällen godkänt stöd till stålföretag som inte tillhör de kategorier som åsyftas i reglerna .
Med omsorg om jämlikhet borde reglerna för statsstöd antingen tillämpas strikt eller ändras , om kommissionen vill godkänna andra stöd än dem som just nu är rättsligt tillåtna .
Slutligen problemet med att EKSG-fördraget löper ut .
Stödsystemet bör finnas kvar efter år 2002 .
På denna punkt är det min uppfattning att endast en förordning från rådet kan ge erforderlig rättslig säkerhet och garantera ett formellt förbud mot alla de stöd som inte täcks av gemenskapens regler .
Av alla dessa skäl har jag röstat för Langenbetänkandet , och jag förväntar mig nu att kommissionen bemöter våra förfrågningar och krav .
( Sammanträdet avbröts kl .
13.05 och återupptogs kl .
15.00 . )
 
Oljebälte vid franska kusten Nästa punkt på föredragningslistan är kommissionens uttalande om oljebältet vid franska kusten .
Härmed överlämnar jag ordet till kommissionens företrädare de Palacio , som får inleda debatten .
Herr talman !
Jag vill börja med att tacka för att parlamentet gett mig möjlighet att tala om den katastrof som inträffat på den franska kusten till följd av förlisningen av oljetankfartyget Erika den 12 december 1999 , något som har lett till att mer än 400 kilometer av kusten har förorenats av den olja som rann ut , att tusentals fåglar har dött , och enormt negativa effekter för miljön och bevarandet av våra hav och hälsosamma kuster som uppfyller de minimikrav som bör kunna ställas i ett välutvecklat samhälle .
Förlisningen av Erika utgör på sätt och vis en antites om det vi alla kämpar för : en hållbar utveckling , en utveckling med respekt för miljön .
Det är ett tydligt exempel på ett brott mot detta sätt att betrakta utveckling och framsteg , ett tydligt exempel på hur det inte får gå till .
Jag skulle kunna lägga ut texten om konkreta fakta som gjorde denna händelse möjlig .
Det kommer jag inte att göra .
Dessa fakta känner vi alla till , och det enda jag vill påpeka är att kommissionen känner samma indignation , inte bara som de som bor vid floden , som är de som i första hand har drabbats av katastrofen på den franska kusten , utan även som alla européer - och inte bara européer - inför en händelse som denna .
Kommissionen visade omedelbart prov på sin solidaritet och har med alla tillgängliga medel försökt stödja bekämpandet av de tragiska följderna av olyckan .
Enligt min uppfattning räcker det inte med att bekämpa följderna , utan det handlar om att komma med lösningar och förslag som gör att man på bästa sätt kan förhindra att dylika händelser upprepas .
Det kan ur miljösynpunkt sägas att vår miljöansvariga kommissionär Wallström omedelbart efter förlisningen bildade en miljökrisgrupp i samarbete med och på begäran av de franska myndigheterna .
Denna grupp startade arbetsgruppen " Havsföroreningar " och ställde de bästa europeiska experterna till de franska myndigheternas förfogande i kampen mot föroreningarna .
Kommissionen medverkade även till att utveckla instrument för bekämpning av föroreningarna på platsen för katastrofen , genom att samordna insatserna från elva av unionens medlemsstater som till platsen skickade mer än 26 kilometer länkar som flyter på vattnet och hindrar oljan från att sprida sig .
Vi anser att denna samordning och resultatet av denna är tecken på framsteg och framgång så tillvida att det verkligen existerar en äkta europeisk solidaritet .
Denna situation är delvis frukten av det arbete som kommissionen bedriver sedan många år tillbaka .
Det arbetet har i synnerhet tagit sig uttryck i upprättandet av ett gemensamt system för insamling av information om alla de stridsmetoder som gemenskapen förfogar över vid den här typen av föroreningar , i tillsättandet av en arbetsgrupp och i den gemensamma finansieringen av projektet för utbildning i och förbättrande av stridstekniken mot föroreningar inom Europeiska unionen .
Förutom lösningar i en nödsituation , är det viktigt att man i längden tillvaratar vår kapacitet att hantera andra liknande katastrofer .
Därför gläds kommissionen över det positiva mottagande som förslaget till beslut om införandet av rättsliga ramar för ett ökat samarbete i bekämpandet av föroreningar till följd av olyckan fick av Europaparlamentet i första behandlingen .
Kommissionen hoppas att de senaste händelserna påskyndar ett slutligt godkännande av denna text i parlamentet och i rådet , och att de nuvarande hindren därmed kommer att undanröjas .
Om vi skall övergå till att tala om transportfrågan , vill jag påstå att förlisningen av Erika på nytt aktualiserar problemet med att förhindra olyckor till havs och rent konkret med säkerheten vid transport , i det här fallet till havs , av förorenat gods .
I den här frågan är det i första hand viktigt att poängtera att Europeiska unionen inte har förhållit sig passiv sedan den omtalade förlisningen av Amoko Cadiz år 1978 , även den utanför den franska kusten .
Kanske bör vi ifrågasätta om man inte borde göra mer , det vill säga om inte vi borde göra mer .
Under de senaste sex åren har ett femtontal förordningar och gemenskapsdirektiv antagits .
Denna lagstiftning är fortfarande ny .
Staterna förfogar i dag över ett rättsligt underlag som gör att de kan ta strid mot bekvämlighetsflagg och mot alla som inte iakttar sina skyldigheter på säkerhetsområdet .
Nu är det upp till medlemsstaterna att visa att det finns en politisk vilja att förse sjöfartsmyndigheterna i respektive stat med de resurser som krävs för att fullföra uppgifter som inspektioner och tillämpning av gemenskapsbestämmelserna , samt en vilja att tillämpa och på lämpligt sätt kräva efterlevnaden av de gemenskapsbestämmelser som redan har antagits .
Kommissionen bör givetvis se till att det sker en enhetlig tillämpning av dessa bestämmelser i samtliga medlemsstater .
Vad beträffar Erikas förlisning har kommissionen redan fått ta del av resultaten från den preliminära undersökning som gjordes av de franska myndigheter om orsakerna bakom olyckan .
Av rapporten framgår hur slarviga - för att använda en eufemism - inspektionerna har varit i det här fallet .
Jag vill påpeka att kommissionen sedan den 21 december 1999 har vänt sig till de italienska myndigheter som är ansvariga för inspektionerna i hamnarna , samt till klassificeringssällskapet RINA , som ansvarar för de senaste klassificeringarna av Erika , för att få en förklaring på hur inspektionerna av Erika gick till .
Faktum är att kommissionen bör ta reda på om de relevanta gemenskapsdirektiven tillämpades på rätt sätt i det här fallet , såväl av de italienska myndigheterna som hamnstat som av sällskapet RINA som klassificeringssällskap .
En sådan undersökning , herr talman , är av största betydelse för att direktiven i framtiden skall kunna förbättras så att vi därigenom också kan förbättra våra insatser .
Hur som helst vill jag meddela parlamentet att en särskild delegation från kommissionen kommer att ge sig av för att granska sällskapet RINA den 28 : e nästa månad och att vi därefter , beroende på vad delegationen kommer fram till , skall vidta lämpliga åtgärder .
När jag säger att vi " skall vidta lämpliga åtgärder " inbegriper jag möjligheten att stryka sällskapet RINA från kommissionens egen lista över kompetenta sällskap .
Dessutom har kommissionen , mina damer och herrar , framfört en liknande begäran till sjöfartsmyndigheten på Malta -Erikas bekvämlighetsflagg - där de hittills , det får jag lov att medge , har varit ytterst samarbetsvilliga .
Utan att på förhand vilja bedöma resultaten av alla undersökningar- hur förlisningen gick till , vilka de yttersta orsakerna var och hur man gick tillväga vid de inspektioner som utfördes , såväl av sällskapet RINA som av de italienska hamnmyndigheterna - så tyder allt på att olyckan med Erika har avslöjat både det ena och det andra som är värt att begrunda och som - enligt min uppfattning - tvingar oss till ett skyndsamt agerande .
Mina damer och herrar , kommissionen höll på att förbereda ett meddelande om säkerheten till sjöss , om säkerheten i hamnarna .
Men det som hänt har tvingat oss att påskynda framläggandet av detta meddelande och i första hand koncentrera oss på transport av farligt och förorenat gods , och då i synnerhet olja , gas och kemikalier .
Detta dokument kommer att åtföljas av en rad lagstiftningsförslag i syfte att stärka sjösäkerheten i gemenskapens farvatten .
Kommissionen räknar med att kunna anta detta innan juni i år , och det innebär att debatterna om de föreslagna åtgärderna , både här i parlamentet och i rådet , kan inledas under andra halvan av år 2000 , under det franska ordförandeskapet .
Vad beträffar innehållet i meddelandet har vi för avsikt att koncentrera oss på följande frågor : I första hand , stärkta kontroller av riskfartyg , oavsett vilket flagg de bär - men det finns statistik som talar för sig själv : av inspektionerna i hamn är felkvoten för fartyg med flagg från en av Europeiska unionens femton medlemsstater cirka 5,9 av 100 utförda inspektioner .
Det internationella genomsnittet ligger på omkring 15,6 för inspektioner som har utförts i europeiska hamnar .
I fallet med fartyg med flagg från Malta - som i Erikas fall - ligger felkvoten på 19,7 och för andra flagg är siffran ännu högre än så .
För att kunna stärka kontrollerna måste vi ändra de gällande direktiven angående klassificeringssällskap , inspektioner av fartygen i hamn och kontrollfrekvensen i förhållande till fartygets ålder och flagg .
När det gäller bilar , måste man som vi alla vet låta besiktiga bilen varje år när de fyra första åren har gått .
Tyvärr är situationen inte den samma för båtar .
Vi förespråkar därför ett liknande förfaringssätt - som å andra sidan har införlivats i de senaste internationella avtalen som ingåtts under IMO : s mantel ( Internationella sjöfartsorganisationen ) genom avtalen SOLAS ( International Convention for the Safety of Life at Sea ) och MARPOL ( en internationell konvention om förhindrande av havsföroreningar från fartyg ) - och se till att detta förfaringssätt blir obligatoriskt .
För det andra bör man främja användningen av miljövänliga oljetankfartyg i de europeiska hamnarna .
Det betyder att de oljetankfartyg som anlöper våra hamnar bör byggas om till oljetankfartyg med dubbelskrov , i stället för att som nu ha ett enkelskrov som innebär att risken för föroreningar är större vid en eventuell olycka .
Den senare typen borde bli föremål för åtgärder för att påskynda ett successivt övergivande av denna , så som sker i Förenta staterna , så att vi undviker den risk vi för närvarande löper : att trafiken med oljetankfartyg som inte kan anlöpa nordamerikanska hamnar omdirigeras till de europeiska hamnarna .
För det tredje , mina damer och herrar , kommer vi i meddelandet att ta upp den komplicerade och känsliga frågan om ansvar och skadeersättning vid en föroreningskatastrof .
Kommissionens avsikt är att ta sig ur denna juridiska härva och lägga fram förslag om att kräva de inblandade parterna på ett större ansvar och dessutom tillsätta nya ansvariga i den kedja där nästan hela ansvaret för närvarande faller på rederiet och fartygsägarna .
Vi har med andra ord för avsikt att införa ett system som gör det möjligt att definiera ägarens eller speditörens ansvar och utkräva detta - om det finns rederier med bekvämlighetsflagg beror det på att det finns fartygsoperatörer som inte fäster något avseende vid kvaliteten på de fartyg de chartrar - samt att öka det antal försäkringar som tecknas av rederierna i förhållande till det totala antalet försäkringar per fartyg .
Kommissionen kommer slutligen att framhärda i sina försök att öka insynen beträffande kvaliteten på de fartyg som trafikerar de europeiska farvattnen .
I det sammanhanget har kommissionen för avsikt att påskynda införandet av systemet Equasix , som bör vara färdigt att tas i bruk i maj i år ; det rör sig helt enkelt om ett system för konkret information i realtid om tillståndet för den internationella flottan med alla dessa båtar .
Programmet håller på att utvecklas i samförstånd med de franska myndigheterna , och innebär att man kan få fram högst konkret fullständig information i realtid om de olika båtarnas tillstånd , för att inte tala om utbildningen av besättningen , som också är en viktig faktor .
Mina damer och herrar , sammanfattningsvis kan jag säga att det inte bara handlar om att diskutera katastrofen med Erika och det som hittills har gjorts , utan även om att dra lärdom så att vi kan undvika en upprepning av katastrofer av det här slaget .
Vi måste garantera en effektiv tillämpning av bestämmelserna för säkerheten till sjöss .
Internationella sjöfartsorganisationen har - som vi alla vet - inte möjlighet att utföra inspektioner eller göra de normer tvingande som antagits av vissa stater där man ofta glömmer sina åtaganden eller inte låtsas om - milt uttryckt - innebörden av de konventioner man har undertecknat .
Dessutom bör vi fortsätta vår strävan efter en ökad konkurrenskraft inom den europeiska rederisektorn , som är en sektor med hög kapacitet och god säkerhet , genom att behålla samma krav som nu , men vi bör också ha förmåga , vad bekvämlighetsflaggen beträffar , att bekämpa det missbruk som uppstår under sådana flagg .
Till slut , mina damer och herrar , gäller det att kämpa mot ett bristande ansvarstagande hos vissa rederier , vissa fartygsoperatörer , vissa stater , vissa sällskap , vissa aktörer på sjötransportens områden som genom sitt bristande ansvarstagande riskerar vår naturliga omgivning och därmed kan förorsaka katastrofer av det slag som olyckligtvis har drabbat den franska kusten på senare tid .
Herr talman !
Jag uttalar mig å PPE-gruppens vägnar , men också i egenskap av förtroendevald från Bretagne som är direkt berörd och chockad av dessa händelser .
Tillsammans med Franoise Grosstête och PPE har vi ingivit ett resolutionsförslag .
I dag har vi ett kompromissförslag framför oss , vilket gläder mig .
Erikas haveri är en europeisk angelägenhet , dels för att det förvanskar och smutsar ned några av Europas vackraste stränder , med mycket allvarliga konsekvenser för turismen , dem som har havet som sin utkomst och de som försvarar miljön , och dels för att detta handlar om regler och kontroller som naturligt sett bör vara europeiska .
En katastrof som denna skulle i princip inte ha kunnat inträffa utanför de amerikanska kusterna .
Varför ?
Därför att amerikanerna har tagit lärdom av Exxon Valdez-katastrofen och därför att de år 1990 utarbetade Oil Pollution Act .
Denna akt utkräver ett större ansvar då den kan göra befraktaren ansvarig , den är dessutom mer tvingande och framför allt bättre kontrollerad genom en rad förordningar och i synnerhet den amerikanska kustbevakningen .
Hade vi haft sådana bestämmelser , jag upprepar detta , hade katastrofen utan tvivel aldrig inträffat .
Därför anser jag att vi måste se över de tillämpliga texterna , och särskilt det protokoll från 1992 som fråntog befraktarna allt ansvar , i det här fallet oljebefraktaren .
Om befraktaren inte är ansvarig blandar han sig givetvis mindre i de kontroller som ligger på oljebolagens ansvar .
Vi måste således se över bestämmelserna , och jag tackar er , fru kommissionär , för att ni pekade på alla de nuvarande bristerna i de europeiska bestämmelserna .
I övrigt krävs det , vilket ni nämnde , framför allt förstärkta kontroller - de kontroller som utförs av den stat under vars flagg fartyget seglar och de som utförs av klassificeringssällskapen .
Ni sade att RINA var ett italienskt klassificeringsregister som har godkänts av kommissionen .
På vilka grunder ges detta godkännande ?
Vilka är garantierna om driftsäkerhet ?
Ni kommer att sända en delegation .
Vi väntar på resultaten med stort intresse .
Man bör också stärka kustmyndigheternas kontroll och kontrollen i europeiska hamnar .
Man skall komma ihåg att det finns en skrivelse från Paris som förutsätter en minimikontroll : en fjärdedel av de båtar som lägger ut från en europeisk hamn måste kontrolleras av det berörda landets kustmyndigheter .
Denna förpliktelse respekteras inte , varken i Frankrike eller i många andra europeiska länder .
Varför ?
Frågan är bara vilka konsekvenser kommissionen redan har tagit eller är beredd att ta ?
Det förefaller också nödvändigt att förstärka den kontroll som befraktaren ansvarar för , i det här fallet oljebolaget .
Om det har ett finansiellt ansvar , kommer denna kontroll utan tvivel att bli bättre .
Till sist krävs det en samordning mellan olika kustmyndigheter för att nå fram till en europeisk gruppering , i likhet med de kustvakter som övervakar Förenta staternas kuster .
För det första skulle jag vilja tacka miljökollegerna i min grupp som tillsammans med sitt transportteam tog tag i detta speciella problem .
Katastrofen är både en transport- och en miljökatastrof och den begränsas inte till ett område .
Så är vi då här igen i detta parlament och diskuterar ännu en sjöfartskatastrof .
Jag skulle kunna rabbla upp en lista på katastrofer som har drabbat denna industri under mina 10 år i parlamentet , men jag har bara tre minuter på mig .
Nu måste det väl vara dags att inte bara medlemsstaterna utan också den där papperstigern som går under namnet Internationella sjöfartsorganisationen och sist men inte minst oljebolagen och tankfartygens ägare tar sitt ansvar och agerar för att stoppa dessa ekologiska och mänskliga tragedier som upprepas år efter år .
Hur många fler Erika måste vi stå ut med innan makterna i fråga ger oss en ordentlig hamnkontroll som gäller inom hela Europeiska unionen och inte bara inom vissa delar av den ?
Hur mycket mera föroreningar måste vi stå ut med innan industrin ger oss tankfartyg med separata tankar och dubbla lastrum ?
Hur många flera sjöfåglar skall dö innan rederierna slutar rengöra sina tankar till havs , vilket orsakar mycket mera föroreningar än någon Erika-katastrof , såsom påpekas i resolutionen ?
Även om jag erkänner att vissa framsteg har gjorts på områden som hamnkontroll och miniminormer för besättningar har vi fortfarande vad vår förre kollega Ken Stewart brukade kalla " skammens skepp " som seglar in och ut på Europeiska unionens farvatten : " dåligt bemannade rosthögar " .
Medlemsstaterna måste handla snabbt och beslutsamt .
Våra regeringar måste ställa upp med de finansiella resurser som fordras för att ge oss en effektiv kontroll och de måste också sluta dra benen efter sig på sjösäkerhetsområdet .
Erika-olyckan har inte tagit några människoliv men den kan ha förstört mångas möjlighet till uppehälle .
Precis som Sea Empress och Braer gjorde .
Det är helt klart att alla tre orsakade ekologiska katastrofer .
Min grupp lider med folket i Bretagne som har fått sin hembygd förstörd av denna katastrof , liksom min grupp led med folket i västra Wales och på Shetlandsöarna vid tidigare olyckor .
Är det inte på tiden att vi slutar uttrycka medlidande och börjar dela ut förelägganden för att bli av med dessa skammens skepp så att vi får säkra hav och inte sitter här igen , senare i år , och diskuterar ett nytt resolutionsförslag när ännu ett bekvämlighetsflaggat tankfartyg tragiskt nog sjunker och spyr ut sin råolja över hela havet .
Tiden för resolutioner är förbi .
Nu krävs handling .
Tyvärr är jag rädd att rådet än en gång kommer att underlåta att göra någonting och att vi i framtiden kommer tillbaka för att diskutera ännu en sjöfarts- och miljökatastrof .
( Applåder ) Herr talman !
Varje gång en sådan här katastrof inträffar säger man att det aldrig får hända igen .
I verkligheten kan vi aldrig sätta stopp för olyckor till havs , men det åligger oss alla att dra lärdom när en sådan här olycka inträffar och använda denna lärdom för att minska riskerna i framtiden .
Erika-olyckan var allvarlig , särskilt för de människor i Bretagne som påverkas närmast , men den var förödande för stora delar av Europas djurliv .
Vissa säger att det var den värsta olycka som någonsin har drabbat fågellivet i denna del av Europa .
Det brittiska Kungliga fågelskyddssällskapet tror att så många som 400 000 fåglar , kanske mestadels alkor , kan ha dött .
De bilder många av oss har sett på oljeindränkta fåglar som avlivas av veterinärpersonal var både sorgliga och tragiska .
Vi vill alla ha högsta möjliga standard på fartyg oberoende av vilken flagg de för .
Vi måste kräva efterlevnad av reglerna och se till att principen om att den som förorenar skall betala tillämpas så att ekonomiska straff och vissa incitament används för att sätta press på både rederier och oljebolag så att en bästa praxis införs .
Jag instämmer i vartenda ord kommissionären sade i sina kommentarer , men frågan är hur lång tid det kommer att ta att tillse att åtgärder genomförs för att ta itu med problemet på det sätt hon föreslår ?
Som politiker måste hon påminna sina tjänstemän om hur svårt det skulle bli om hon skulle behöva komma tillbaka till detta parlament om ett år om en liknande , precis lika förödande olycka skulle inträffa , och vissa av de åtgärder hon föreslår i dag fortfarande bara vore vackra ord som hon inte hade haft möjlighet att omsätta i verklighet .
Tanken på att en olycka av detta slag kan inträffa inom en nära framtid bör bidra till att skärpa hennes och hennes tjänstemäns sinnen på ett fantastiskt sätt .
Herr talman , fru kommissionär !
Jag har tagit med en liten present till er : det är en oljekoka som en invånare på ön Noirmoutier har skickat till mig , och hon skriver följande : " varje gång det är flod täcks stranden av tung olja som läckt från Erika .
Varje gång det är flod tar frivilliga , militärer och brandmän fram enorma kokor av denna svarta klibbiga och tjocka tjära .
När blir det rent igen , när blir det ett slut på denna ödesdigra olycka ? "
Ja Erikas haveri , liksom den ryska båtens haveri i Turkiet för övrigt , kan inte accepteras eller tolereras med tanke på att den tekniska utvecklingen står på sin höjdpunkt .
Det är dessutom oacceptabelt om man betänker att olyckan inträffade 20 år efter Amoko Cadiz-katastrofen , när man redan har sagt och flera gånger upprepat : " aldrig mer ! "
Det är självklart politikernas , och därmed vårt ansvar att garantera säkerheten vid transporter till havs .
Vi måste verkligen försäkra medborgarna att en liknande olycka aldrig mer kommer att inträffa .
Men vi blir något frustrerade när vi lyssnar till er , fru kommissionär , för de som redan har ägnat sig åt den här typen av frågor vet att kommissionen och parlamentet förberedde , jag tror det var 1992 , en mycket intressant text , som redan då innehöll alla de förslag som finns i dagens resolution från utskottet för regionalpolitik , transport och turism .
Det måste upprepas och upprepas igen : Erika var en katastrof för mycket .
Därför är det brådskande att Europeiska unionen inleder en genomgripande revidering av direktiven om transporter till havs , för att göra dem mer tvingande samt upprättar en klar och detaljerad ansvarsordning för lastens ägare .
Man bör t.ex. känna till att såväl Shell som British Petroleum vägrade att använda Erika för sina oljetransporter .
Varför medger man inte under dessa omständigheter att befraktaren , Total , har ett ansvar ?
I era förslag bör ni även kräva dubbla fartygsskrov och att förbudet mot tankrengöring till havs verkligen respekteras .
Man måste inrätta en europeisk inspektörskår , så att de verkligen och effektivt kan kontrollera båtarnas skick .
Det är för övrigt lika brådskande att Europeiska unionen åtar sig att reformera Internationella sjöfartsorganisationen ( IMO ) .
För vad tjänar det till att utarbeta bindande direktiv , om sedan flertalet båtar gör vad de vill när de väl är ute till havs ?
Till sist , mina damer och herrar , vill jag skänka en öm tanke till alla frivilliga , natur- och fågelvänner , som spontant och generöst har anmält sig för att rädda oljeindränkta fåglar , genom att organisera en räddning med de medel som står till förfogande .
Jag kan intyga att det är ett anmärkningsvärt arbete .
Ni känner utan tvivel till att omkring 200 000 fåglar kommer att gå under i detta oljebälte , som är en oerhörd miljökatastrof och som praktiskt taget saknar tidigare motsvarighet .
Ni vet också hur svårt det är i dag att bevara djurarter och hur svårt det är att bevara naturområden .
På den punkten , fru kommissionär , sade ni ingenting , dvs. hur kommissionen avser att bidra till återställandet av naturen och livsmiljöerna .
Än en gång kommer ingen ansvarig att utpekas klart och tydligt .
I väntan på det är det alltid naturen som tar stryk .
Herr talman !
Min grupp begärde denna debatt för att ge parlamentet tillfälle att uttrycka sin solidaritet med de personer som är direkt berörda av miljökatastrofen , såväl i sin ekonomiska verksamhet som sina känslomässiga relationer med naturen .
Tillåt mig att välkomna talesmannen för kollektivet " Oljebältet " , bestående av medborgare från departementet Morbihan ; Javette-Le Besque , som har tagit plats på åhörarläktaren .
Att uttrycka sin solidaritet , det har många frivilliga från Frankrike och olika europeiska länder gjort genom att ge en viktig hjälpande hand till de drabbade .
Att uttrycka vår , Europaparlamentets solidaritet , det är i första hand att agera för att omedelbart få fram ett katastrofstöd till de familjer som drabbats av oljebältet .
Det innebär också att kräva en kvalitativ förstärkning av europeiska och internationella regler och säkerhetsnormer för transporter till havs , med tätare kontroller och mycket mer avskräckande sanktioner gentemot dem som bryter mot reglerna .
Våra förslag avser bl.a. oljetankrarnas ålder .
Bland dem som kontrollerades och bedömdes som bristfälliga förra året , var 15 av dem 20 år eller äldre , vissa mer än 30 och t.o.m. ännu äldre .
Det kan inte längre tolereras .
Vidare bekvämlighetsflaggade fartyg .
Enligt Internationella transportfederationen seglade 40 procent av de fartyg som havererade 1998 under bekvämlighetsflagg , en symbol för vinst och utnyttjande av människor till förfång för säkerheten .
Det kan inte längre tolereras .
Slutligen bristen på öppenhet .
Man gör allt för att mörklägga kedjan av ansvariga , ägarnas identitet och de verkliga beslutsfattarna .
Det kan inte längre tolereras .
I alla dessa avseenden måste vi utverka verkliga och betydelsefulla förändringar , bl.a. en tidsfrist för inrättandet av nya normer som dubbla fartygsskrov .
De som inte uppfyller kraven skall inte få lägga ut från hamnarna eller kryssa på medlemsstaternas vatten .
Vi måste också uppnå ytterst strikta regler när det gäller utfärdande av sjövärdighetscertifikat och bedömningen av fartygens skick och underhåll .
Vi måste slutligen se till att alla som bär ansvaret för en katastrof också bidrar till reparationerna .
I det här fallet tänker jag på gruppen Total-Fina .
Herr talman !
Denna strategi kan Europeiska unionen utveckla visavi Internationella sjöfartsorganisationen .
Då kommer vi att ha visat allmänheten att vi gör någon nytta , för den här gången väntar man sig tydlig och konkret handling .
Herr talman , fru kommissionär !
I egenskap av förtroendevald från den franska atlantkusten , från Vendée , vill jag först och främst uttrycka den upprördhet som offren för Erikas oljebälte känner inför katastrofen , en katastrof som har förorsakats av - inte en naturkatastrof som de orkaner vi nyligen drabbades av - utan av en brottslig handling .
I det akuta läget och inför en stor prövning , uttrycktes en fantastisk solidaritet : en lokal solidaritet , en nationell solidaritet , en mellanstatlig solidaritet .
Förväntningarna hos de drabbade befolkningarna , de som har förlorat allt - särskilt de som är yrkesmässigt beroende av havet och turismen - de vilkas verksamhet är ruinerad för flera år framöver , är inte bara att förorenarna skall betala för de skador de har åsamkat , utan också att man gör allt för att deras olycka skall hjälpa andra i framtiden och förhindra att liknande brott begås igen .
Vi betalar givetvis priset för våra försummelser .
Staterna gjorde nämligen bedömningen - med gemenskapens välsignelse - att det inte längre var lönsamt att ha en egen handelsflotta och lät därmed ett stort kunnande i skeppsbyggnad försvinna .
Därför kan vi inte längre spåra fartygens ursprung och därför får vi se riktiga vrak segla på våra farvatten under bekvämlighetsflagg , till förmån för de multinationella bolagens kortsiktiga intressen .
Vi måste verkligen sätta stopp för denna ström av oansvarighet , oansvariga befraktare , skeppsredare som är omöjliga att hitta och eftergivna certifieringssällskap .
Dagens läge är mycket förvirrat .
Dessa frågor bör självklart hanteras på internationell nivå , men IMO : s nuvarande internationella regler är otillräckliga och alltför släpphänta .
Varken medlemsländerna eller gemenskapen har varit påstridiga och försökt få till stånd striktare regler , trots tidigare inträffade katastrofer .
Visserligen existerar Internationella fonden mot oljeföroreningar ( FIPOL ) , men den sprider ut ansvaret och har alltför begränsade ramar , som därför måste ses över .
Man bör absolut se över frågan om bekvämlighetsflagg inom ramen för IMO .
Det är medlemsstaternas och gemenskapens sak att vidta erforderliga åtgärder för det ändamålet .
Jag vill erinra om att Erika bekvämlighetsflaggades av en stat som har ansökt om medlemskap i unionen .
Vi har också gemenskapens direktiv , men de tillämpas i ringa utsträckning eller inte alls , på grund av att de nationella kontrollanterna är alltför få .
Vi måste snarast åtgärda den bristen .
Ett direktiv om säkerhet till havs har förberetts under många år , men arbetet framskrider mycket långsamt .
På den punkten visar kommissionen en tröghet som inte kan tillåtas och en oförmåga som inte kan accepteras .
Presentationen av kommissionens meddelande om denna centrala fråga skjuts ständigt upp och är nu planerad till juli , men den bör absolut tidigareläggas .
Vad gäller de konkreta bestämmelserna måste de vara särskilt tydliga och strikta .
Jag vill nämna tre som vår grupp prioriterar .
För det första måste tankerägarnas ansvar klart och tydligt fastställas , och de som faller offer för en förorening måste utan tvekan kunna ställa dem till svars .
Det bästa sättet att förebygga olyckor inför framtiden , är att befraktarna kan vara förvissade om att de kommer att straffas hårt , civilrättsligt , straffrättsligt och finansiellt , om de inte är ytterst vaksamma beträffande säkerheten på de fartyg de väljer ut .
För det andra måste kravet på dubbla fartygsskrov för oljetankrar som får segla på gemenskapens farvatten införas så snart som möjligt , och inte uppskjutas på obestämd tid .
För det tredje måste man snarast fastställa en strikt begränsning av åldern på de fartyg som tillåts frekventera gemenskapens farvatten .
Maximiåldern skulle kunna vara 15 år .
Lyckas man inte uppnå en tillräckligt tydlig , strikt och rigorös ram på gemenskapsnivå , bör de medlemsstater som för egen del vill införa striktare bestämmelser tillåtas att göra det för att skydda sin befolkning och sitt territorium , på samma sätt som Förenta staterna tog lärdom av Exxon Valdez-katastrofen genom att kräva dubbla fartygsskrov och förbjuda alla fartyg som är äldre än 20 år att segla på deras farvatten .
Förenta staterna skulle således ha vägrat Erika tillträde till sina farvatten .
Om gemenskapen hade gjort detsamma hade en oerhörd katastrof kunnat undvikas .
Herr talman , fru kommissionär !
Låt oss denna gång verkligen ta lärdom , även när massmedias och parlamentsledamöternas känslor har lagt sig .
Herr talman !
Torrey Canyon , Olympic Bravery , Haven , Amoko Cadiz , Gino , Tanio ; detta är en rad namn som är förknippade med dystra minnen .
Och nu Erika .
Vems tur är det sedan ? 21 år efter Amoko Cadiz får vi för femtielfte gången se ett oljebälte , det sjunde sedan 1967 och beviset för alla efterföljande regeringars oansvarighet .
Västra Atlanten får än en gång betala ett högt pris för deras oförmåga att reagera , för att de kapitulerar inför de multinationella bolagen .
Det är svårt att förstå varför fransmännen och européerna tillåter det som amerikanerna förbjuder , och varför Europa , som normalt sett är så snabbt på att lagstifta i miljöfrågor , inte har gjort något för säkerheten till havs .
Resultatet ser vi i dag .
Erika , ett fartyg som seglade under maltesisk flagg , ett flytande vrak som klassas som en av de farligaste oljetankrarna , har smutsat ned våra kuster längs en drygt 400 km lång sträcka , vilket är en långt mer allvarlig förorening än den som Amoko Cadiz förorsakade .
Som förtroendevald från Loire-Atlantique kan jag tyvärr intyga det .
Dessa upprepade katastrofer hänger på inte på något sätt samman med naturens krafter , det finns inget ödesbestämt över dem .
De är en konsekvens av människors inkonsekvens .
Detta är en riktig miljökatastrof .
Endast de som inte har varit där och sett den hårda verkligheten kan betvivla det .
Det är också en ekonomisk katastrof för alla dem som lever av havet och turismen ; fiskare , ostronodlare , musselodlare , salinarbetare , handlare , osv .
Svepeskålen Erika måste bli den sista i raden .
Vi måste först och främst göra allt för att bringa klarhet i haveriet .
Varför inte utse en parlamentarisk undersökningskommitté eller låta parlamentsledamöter delta i den delegation som kommissionen aviserade för en stund sedan ?
Sedan måste vi snarast anta lagar som fordrar grundligare kunskaper om det transporterade godsets egenskaper .
Enligt experterna skulle oljan från Erika ha sjunkit till bottnen och aldrig ha nått kusterna .
Men vi vet vad som hände .
Det krävs vidare att man inför en tillförlitlig teknisk kontroll , i likhet med Frankrikes obligatoriska tekniska kontroll av fartyg som är äldre än fem år .
Det krävs bestämmelser för användningen av bekvämlighetsflagg , krav på dubbla fartygsskrov för transporter av förorenande och farliga ämnen och en utveckling av tekniken för att hantera och samla upp oljeutsläpp .
Det är enligt min mening ett minimum på tröskeln till det tredje årtusendet .
De fartyg som inte uppfyller kraven måste nekas tillträde till europeiska farvatten ; förorenarnas , skeppsredarnas och befraktarnas ansvar måste fastställas enligt principen " den som förorenar skall betala " ; övervakningen på haven måste förstärkas för att förhindra tankrengöring ; en seriös och tillförlitlig kontroll av fartygstankrarna måste införas ; en konsekvent budgetpost för " naturkatastrofer " måste återupprättas för medlemsländerna , och i väntan på det bör man uppbåda ett exceptionellt gemenskapsstöd och se till att medel ur strukturfonderna kan anslås till de katastrofdrabbade departementen .
Å EDD-gruppens vägnar har jag också ingivit en resolution i den frågan .
Herr talman !
Under de senaste åren har det över hela världen förekommit upprepade svåra katastrofer med tankfartyg , utan att några nämnvärda eller effektiva motåtgärder har vidtagits .
Denna gång är det särskilt illa , inte minst därför att det har drabbat en stor europeisk stat , en händelse som kan upprepas när som helst .
För att minska dessa risker behöver vi snarast ett direktiv .
De 15 räcker uppenbarligen inte .
Dessa garanterar - utan anspråk på att vara fullständiga - minst 3 punkter : Inget skrotfärdigt tank- eller fraktfartyg får någonsin mer anlöpa en hamn i Europeiska unionen .
Alla inblandade , inklusive den som beordrat transporten , är ansvariga för följdskadorna , och tillräckliga försäkringar måste tecknas av dessa inblandade .
Endast på så sätt kan de drabbade ha en chans att få sina skadeersättningsanspråk tillgodosedda .
Men vi måste vara klara över att det långsiktiga målet måste sättas mycket högre .
Det betyder att vi behöver en verklig kostnadsuppskattning för vårt hela energiförsörjningssystem .
Herr talman !
Skulle jag kunna få börja med att rikta ett stort tack till kommissionär Palacio för det klara , adekvata och även mycket rakryggade svaret .
Tusen tack för detta .
Det innebär också att jag i varje fall har stor respekt för det briefing-PM som hon skickade den 10 januari , men också för de åtgärdspunkter som hon tillkännagav i dag .
Katastrofen med Erika visar att när övergripande trafik- och transportbestämmelser saknas på internationell och europeisk nivå så är det naturen och miljön som drar det kortaste strået .
Den skada som har uppstått , även på det ekologiska området , går inte att uttrycka i pengar .
Det är anledningen till denna gemensamma debatt med kollegerna från transport och miljö .
Under julferien när de nederländska medierna uppmärksammade katastrofen med Erika gick jag ut på Internet för att se vilka åtgärder det nu egentligen var som skulle vidtas , i synnerhet efter det att premiärminister Jospin hade sagt att Europa måste göra mer .
Vad jag förstod av detta var att det egentligen finns tillräcklig lagstiftning , men att problemet är att det inte sker några kontroller .
Jag skulle här vilja uppmärksamma ett par punkter , som även kommissionären nämnt i förbigående .
Först och främst port-state control , de 25 procent av alla fartyg som måste kontrolleras .
Jag tror att dessa 25 procent inte bara måste upprätthållas , utan att man därefter också måste sörja för att det görs fler kontroller ; dessa 25 procent måste således höjas .
När ett skepp inte längre får segla måste inte bara sakförhållandena kontrolleras , utan det måste också inrättas ett rättsligt system där man säger : det är klokast att ni inte går ut till havs mer eller det får ni inte göra längre .
Men något sådant finns inte .
Herr talman !
På den punkten skulle jag gärna se att det hände något .
Slutligen något om de tekniska krav som ställs på fartyg ; mina kolleger talade nyss om att det i Förenta staterna sedan 1999 i varje fall måste finnas dubbla kölar .
Jag anser att vi måste gå längre på den punkten , och jag anser också att Marpol-fördraget , som träder i kraft 2001 , måste ses över ordentligt .
Herr talman !
Sedan måste man också kritiskt se över anslutningsförhandlingarna med Malta , och jag vill framföra mitt tack och min beundran till de många icke-statliga organisationer som i varje fall har tagit upp händerna ur byxfickorna för att rädda djur .
Herr talman !
Vi har redan ofta fört denna diskussion .
Vi har hittills inte uppnått någonting , och vi har inte kunnat enas här i Europeiska unionen .
Därför tror jag att det bara är meningsfullt med dagens debatt om det som vi alla säger i dag , och det som ni , fru kommissionär , här har tillkännagett , faktiskt utmynnar i en lagstiftning , dvs. om ni säger till alla era regeringschefer och era ministrar : Detta måste ni genomdriva i ministerrådet .
Låt mig på förhand säga att vi talar om en miljökatastrof , som också har ekonomiska effekter och hotar existenser .
Vad måste vi nu göra ?
Jag vill ju alls inte gå tillbaka till det förflutna .
Jag vill se framåt .
Vad skall vi göra nu ?
Jag vill säga något om vad vi måste göra .
Naturligtvis behöver vi fartyg med dubbelt skrov .
Det är klart , men detta är något som bara kommer att få effekt på medellång och lång sikt .
Vad behöver vi då genast ?
Vi behöver en teknisk kontroll av fartygen , nämligen en bindande teknisk kontroll av fartygen vartannat år , och utan detta certifikat får inget fartyg framföras .
Det behöver vi på europeisk nivå , och det behöver vi internationellt , som en teknisk övervakningsinstans , som en teknisk besiktning av fordon , vilken i Tyskland måste göras vartannat år .
Om man inte har något besiktningsinstrument , får man inte köra fordonet .
Det behöver vi för fartyg .
För det tredje behöver vi en kontroll av dessa certifikat och ett försäkringsbevis i hamnarna , och detta i alla Europeiska unionens hamnar .
Om detta certifikat och försäkringsbevis saknas , beläggs fartyget med kvarstad och får trots alla hamnavgifter inte lämna hamnen .
Där måste vi vara ense , i alla hamnar i Europeiska unionen , från Marseille via Rotterdam till Wilhelmshaven , Cuxhaven och var än fartygen anlöper .
För det fjärde måste det finnas ett ansvar hos fartygsägaren , och inte bara skrattretande 12 miljoner dollar , utan minst 400 miljoner dollar , vilket han måste styrka med hjälp av försäkringsbevis .
Då måste det finnas ett ansvar hos det land , under vars flagga fartyget seglar .
Vi behöver den säkerheten att det land , under vars flagga fartyget seglar , i tveksamma fall övertar ansvaret .
Det blir en underbar kontroll !
Jag kan garantera att de länder som utdelar flaggorna då också kommer att se till att de inte måste bära ansvaret .
Vi behöver för det femte den garantin att detta krävs för alla fartyg i Europeiska unionens hamnar och farvatten , för övrigt också i kandidatländernas .
Det betyder att de krav som jag har nämnt gäller för alla farvatten .
Slutligen behöver vi det allra viktigaste : Vi behöver ha ett bra minne , ty vi kommer här under den närmaste tiden att oftare tala om lagstiftning .
Vi kommer oftare att tala om miljönormer .
Då vill jag inte att någon kommer och säger : Dessa krav leder till att vi förlorar arbetstillfällen i hamnarna .
Fackföreningarna kommer , industrin kommer .
Vi behöver ett bra minne , kära kolleger .
Här tittar jag på många av er , som hittills inte har gått i bräschen för miljörörelsen .
Gå hem och säg : De normerna har vi hittills inte bekymrat oss om .
Vi behöver ett bra minne när det gäller vad som krävs i hamnarna .
Vi behöver ett bra minne , när vi säger : Vi är ense vad beträffar hamnavgifter och hamnbestämmelser , och vi spelar inte ut den ena mot den andra i Europeiska unionen .
Om vi klarar av det , så kommer vi kanske om ett par år att ligga bättre till !
Herr talman !
Roth-Behrendt uttryckte väldigt mycket av mina tankar .
Vi har nu fått en perfekt uppräkning av olika åtgärder .
Men hur använder vi det krismedvetande som denna ekologiska katastrof har lett till ?
Jag jämför med när en tidigare generation införde plimsollmärket , en märkning som infördes för att undvika försäkringsbedrägerier med undermåliga fartyg .
Var har vi samma krismedvetande som generationerna före oss hade ?
Jag anser att det vi skall gå in för är den certifiering som Roth-Behrendt talar om , den märkning med gröna märken på tankfartyg som vissa hamnar i Europa har fört på tal .
Vi måste dessutom kritiskt granska klassificeringssällskapen .
Jag tycker inte att vi kan acceptera deras förfarande .
Vi behöver oberoende förfaranden och förfaranden med insyn .
Slutligen vill jag säga att när mitt land ger miljöstöd till redare som vill förbättra miljökvaliteten , så finns det enheter inom kommissionen som betraktar detta som förbjudet varvsstöd .
Den ena handen inom kommissionen vet inte vad den andra gör .
Det är inget acceptabelt förfarande att man inte får göra miljöförbättrande åtgärder , som är i enlighet med kommissionens riktlinjer , eftersom dessa anses utgöra förbjudet varvsstöd .
Herr talman !
Vi kommer att rösta för resolutionen från GUE / NGL-gruppen , eftersom den pekar ut Total-Fina som ansvarig för denna miljökatastrof , och eftersom jag skriver under på förslaget att förbjuda bekvämlighetsflagg och bruket av föråldrade båtar , och att införa ett krav på dubbla fartygsskrov för oljetankrar .
Jag vill bara tillägga att det minsta man kan begära är att Total betalar alla kostnader för de skador som oljebältet direkt och indirekt har förorsakat .
Hur skall man kunna förhindra att liknande katastrofer inträffar igen om man inte vidtar ytterst stränga åtgärder gentemot de stora oljetrusterna , och även andra , som för att kamma in ytterligare vinster tar risken att göra vår planet obeboelig ?
Hur är det möjligt att inte uppröras över att en bank vägrar lämna ut namnet på Erikas ägare genom att hänvisa till banksekretessen , och att ingen regering reagerar på det ?
Det egentliga problemet är att alla regeringar , liksom alla EU-institutioner , ger stora truster som Total-Fina och dess likar rätten att maximera vinsterna till nackdel för såväl sina anställda som miljön .
Man tillerkänner företag och banker rätten att hemlighålla sina affärer , även om denna sekretess skyddar rent kriminella handlingar .
Under dessa omständigheter kommer även de allra bästa resolutioner att förbli bevisningsfel , som inte kan förhindra att de stora trusterna åsamkar skador .
Herr talman , kära kolleger !
Jag anser att vi bör skärpa föreskrifterna om hamnstatskontrollen och om organisationerna som utför inspektionerna .
Men vi måste också se på fakta .
Fartyget Erika hade undersökts fyra gånger under de senaste två åren .
Det är inte antalet undersökningar som är avgörande , utan det är snarare så att intensiteten i kontrollerna måste garanteras .
Under diskussionerna de senaste veckorna har jag hört sägas att medlemsstaterna inte har tillräckligt med pengar för att genomföra kontrollerna !
Det kan jag inte acceptera .
Om medlemsstaterna gemensamt med oss beslutar att 25 procent av fartygen skall kontrolleras på grundval av hamnstatskontrollen , då måste de också ställa personal till förfogande !
Då måste kontrollerna också genomföras så att inspektören inte bara går ombord och tittar efter om det möjligen saknas en brandsläckare , utan då måste det göras materialprovningar , ty detta fartyg har uppenbarligen brutits isär på grund av materialutmattning .
Det kan man bara fastställa med hjälp av intensiva kontroller .
Det bör vara vårt mål att se till att hamnstatskontrollerna inte är ytliga , utan att man inkluderar materialet .
För det andra håller jag också med om kommissionärens antydningar och vill uppmuntra henne att fortsätta på detta vis .
Om det skulle visa sig att en eller flera organisationer som utövar tillsynen har avgett vänskapsutlåtanden , då skall de strykas från listan med tillåtna organisationer !
Det är det enda sättet att avskräcka organisationerna från att också avge vänskapsutlåtanden .
Kära kollega Roth-Behrendt , vi har en teknisk övervakningsinstans för fartyg .
Organisationerna som skall utföra inspektionerna är den tekniska övervakningsinstansen för fartyg !
Det finns också bra organisationer .
Du känner till några bra organisationer , våra franska kolleger känner till några bra organisationer , men vi måste se noga efter vilka organisationer som inte uppfyller villkoren , och dessa måste strykas från listan .
En sista punkt : Vi bör entydigt säga till Malta att om Malta vill bli medlem av denna gemenskap så måste det fram till anslutningen tillämpa en standard vid registreringen och vid flaggstatskontrollen som verkligen motsvarar våra anspråk , ty miljön är gemensam för oss , och ingenting man kan dela upp !
( Applåder ) Herr talman , fru kommissionär !
Erika sjönk rakt framför mitt hem .
Hon ligger fortfarande där med 20 000 ton i sidorna , och man vet ännu inte vart dessa ton kommer att ta vägen .
Hon hade kunnat sjunka någon annanstans .
Men av en slump sjönk hon just där , och det Bretagne som jag kommer ifrån skall inte behöva ursäkta sig för att det är en halvö , för Bretagne får ofta uthärda skeppsbrott .
Jag tänker framför allt på de 26 indiska sjömän som man inte talar om och som inte räddades .
Människor hade kunnat dödats i den här katastrofen , och säkerhet till havs handlar främst om människoliv .
I dag är dessa sjömän ett avlägset minne .
Det är ett mirakel om de har räddats .
Så kommer man att börja om på nytt precis som för 20 år sedan med Amoco , ett hugg på nordkusten , ett hugg på sydkusten , ett hugg på västkusten .
Och det skulle kunna fortsätta på det viset .
Fru kommissionär !
Eftersom det är mycket ont om tid skulle jag bara vilja räkna upp de sju punkter som vi anser att det är ytterst viktigt att arbeta på , och ni har säkerligen nämnt några av dem : dubbla fartygsskrov så snart som möjligt på våra farvatten och en så strikt statlig kontroll som möjligt i hamnarna .
Det krävs framför allt att klassificeringssällskapen är förpliktade att offentliggöra sina rapporter , eftersom de inte är kända .
Vidare att de femton medlemsstaterna harmoniserar påföljderna - de får inte skilja sig åt , utan måste vara desamma överallt .
Man måste skärpa bestämmelserna om bekvämlighetsflagg , inte för att de nödvändigtvis är sämre båtar , utan för att det finns många dåliga båtar som seglar under bekvämlighetsflagg ; förbättra informationen om samtliga fartyg i världen , vilket visserligen redan är planerat , och att ringa in och skärpa ansvaret .
I det avseendet skulle jag vilja veta vem som äger Erika , för begreppet juridisk person i vår rätt är en sak , men det finns alltid fysiska personer bakom - var är de , Erikas ägare ?
Kanske i vackra villor vid vackra stränder för att sola sig .
Vi skulle gärna se deras namn och deras ansikten .
Och slutligen en förbättring av utbildningen för fartygsbesättningar .
I vårt samhälle finns det ingenting som en nollrisk , men vi kan åtminstone vara så försiktiga som möjligt .
Herr talman !
Jag välkomnar kommissionärens uttalande .
Eftersom jag själv har tillbringat lång tid till sjöss är jag väl medveten om havets makt och destruktiva kraft som gör ändamålsenlig utformning och underhåll av skepp och båtar avgörande .
Jag skulle vilja uttrycka mitt deltagande med alla dem som handskas med konsekvenserna av att oljetankern Erika förliste och sjönk .
Detta har varit en miljökatastrof liksom ett djupt beklagligt resursslöseri .
Man bör notera att oljeindustrin , genom de internationella oljeskadefonderna , betraktar sig som ansvarig för över 90 procent av den beräknade kostnaden för denna olycka , eller cirka 170 miljoner dollar , enligt konventionen från 1969 och 1992 års protokoll .
Detta tycker jag tyder på att vi också bör uppmana fartygens ägare , den stat vars flagg man för och kontrollmyndigheterna att ta sin del av ansvaret .
Låt oss emellertid , innan vi rusar åstad med en hel räcka nya åtgärder och regler , noggrant titta på gällande bestämmelser så att vi är säkra på att de tillämpas på rätt sätt .
Det är bättre att följa uppmaningar att modifiera och förbättra gällande lagstiftning än att inlåta sig på nya förslag .
I detta sammanhang stöder jag kraven på att utöka hamnkontrollen för att tillse att en total och effektiv kontroll görs .
Jag stöder krav på att tillse att klassificeringssällskapen på ett effektivt sätt övervakar fartygens strukturella skick och hålls ansvariga för sina handlingar .
Krav på förbättringar av skrovkonstruktionens utformning , speciellt fartyg med dubbla skrov , är förnuftiga men tar tid att genomföra i hela flottan .
Det finns inget som kan ersätta rigorösa regelbundna kontroller .
Herr talman !
Jag vill framföra ett tack till mina socialistiska kolleger , i synnerhet till dem från utskottet för regionalpolitik , transport och turism samt utskottet för miljö , folkhälsa och konsumentfrågor , för att de inte har glömt att denna olycka även påverkar fiskerisektorn .
Förutom skadorna på miljön , skadorna på ekosystemet som inte går att reparera och förlusterna för turistsektorn , innebär oljebältena ett dråpslag för fisket , för bevarandet av resurserna i havsmiljön , och det kommer att ta många år att återställa den förstörda kusten .
Det är ingen tillfällighet , fru kommissionär , att de drabbade områdena alltid är europeiska regioner med en försenad utveckling , de regioner som hankar sig fram med hjälp av en kombination av turism och fiske , och där det i de flesta fall saknas andra resurser .
Det är även dessa regioner , fru kommissionär , som under hela året får stå ut med vissa redares oförskämda agerande då de rengör botten på sina fartyg utanför kusten , utom all kontroll .
Jag kommer själv från Galicien , en region som tidigare har drabbats av liknande olyckor .
Bretagne och Galicien , två europeiska ändpunkter , blir ständigt offer för det bristande ansvarstagandet hos dem som väljer att bryta mot säkerhetsbestämmelserna och transportera råolja i fartyg som i sig utgör potentiella oljebälten .
Därför anser jag att det är nödvändigt att agera i två olika avseenden .
För det första genom att vi ber att kommissionen , inom ramen för det planerade stödet till fiskerisektorn , vidtar särskilda åtgärder för att mildra effekterna av denna katastrof för den produktiva sektorn i de drabbade regionerna , och att vi dessutom ber kommissionen av sig själv och de internationella organen kräva en striktare kontroll av fartyg med bekvämlighetsflagg .
Därför bör man under den pågående förhandlingsprocessen om Maltas anslutning till Europeiska unionen passa på att kräva att Malta utövar en sträng kontroll av oljetankfartyg under deras flagg .
För det andra måste vi agera förebyggande .
Portugal är ett land där man tydligt visat hur känslig man är för frågor med anknytning till havet .
Jag skulle vilja uppmana det portugisiska ordförandeskapet att undersöka möjligheten att införa en övergripande strategi för att förebygga olyckor till sjöss på europeisk nivå , genom att man sammanför all de medel som står till vårt förfogande - tekniska , strukturella och socioekonomiska sådana - för att undvika en upprepning av en katastrof som denna i framtiden .
Slutligen , herr talman , vill jag lyfta fram det arbete som har utförts av frivilliga och av de lokala myndigheterna , som påminner mig om gamla tider då jag - som borgmästarinna - fick uppleva liknande situationer .
Vi måste tacka alla dem som i ett sådant utsatt läge med knappa resurser har visat mod i kampen mot de allvarliga konsekvenserna av denna katastrof för kustregionerna , ekosystemet till sjöss och Europas fiskeresurser .
Herr talman !
I egenskap av ordförande för utskottet för regionalpolitik och transport skulle jag vilja gratulera kommissionen , och speciellt kommissionsledamoten Loyola de Palacio , till deras sätt att hantera denna fråga , som har väckt så starka reaktioner i hela Europa .
Vi i transportutskottet är beredda att diskutera kommissionens meddelande om säkerhet till havs , och vi är naturligtvis också beredda att senare diskutera vilka konsekvenser detta meddelande får i rättsligt avseende .
Sedan skulle jag vilja göra några påpekanden : För det första ; det är med all rätt som kommissionen i sin undersökning framför allt söker utkräva ansvar av det italienska fartygsinspektionsbolaget RINA , eftersom vi måste ta reda på om gemenskapsrätten har tillämpats .
Detta bör vara utgångspunkten för våra ansträngningar .
För det andra ; förutom redarnas ansvar är det lämpligt att vi i sådana fall även beaktar befraktarnas ansvar , det gäller t.ex. oljebolagen som också bär ansvar för ekologiska katastrofer som i det här fallet , men som också måste ta sitt ansvar för att återställa det som skadats .
Reaktionen på den ekologiska katastrofen är verkligen befogad .
Men detta får inte leda till att vi skuldbelägger all handelssjöfart , som ju är en mycket viktig bransch för ekonomin , eftersom den svarar för ungefär 1 / 3 av transporterna , och därför bör våra reaktioner vara måttfulla , stränga men också korrekta .
Jag motsätter mig inte alls att man överväger en skärpning av gemenskapsrätten men , såsom även andra kolleger har framhållit , vi bör utgå från tillämpningen , för det finns redan ett regelverk - och det får vi inte glömma - på Europeiska unionens nivå .
Detta regelverk är ganska avancerat - åtminstone om man jämför det med situationen på global nivå - och följaktligen är medlemsstaterna , under kommissionens överinseende , skyldiga att verkligen börja tillämpa gemenskapsrätten .
Herr talman !
Jag tror att man bara kan välkomna kommissionärens sakliga och nyktra konstateranden , ty hon har inte gjort det som andra gör , nämligen att förfalla till kollektivt hycklande .
Katastrofen med Erika var inte överraskande .
Jag vet inte hur många de är , men en stor mängd fartyg som praktiskt taget utgör flytande tidsinställda bomber far varje dag i europeiska farvatten , och en sådan katastrof kan såvitt vi ser det också upprepas när som helst .
Detta har vi känt till i mer än tio år i detta parlament - det kom då ett meddelande från kommissionen , och ett betänkande från vår kollega Ken Stewart , där alla områden redan nämndes , där man måste utfärda lagbestämmelser .
Och här handlar det om fartygen , tekniken och utrustningen ; det handlar om hamnarna , hur de organiseras och vad som krävs där , och det handlar naturligtvis också om de bra manskapen .
Vi vet mycket väl varifrån motståndet kom i samband med varje enskild laglig åtgärd under de senaste åren .
Motståndet kom alltid från medlemsstaterna , från ministerrådet , där man envist brottades om varje småsak för att uppnå ett litet framsteg .
Om vi å ena sidan begär av varje medborgare som har ett personfordon att han själv måste vara frisk och se till att han har ordentliga personliga förutsättningar , och han å andra sidan måste låta göra en regelbunden besiktning av sitt personfordon , måste detta också vara möjligt för fartyg .
Kontroll är nyckelordet i denna fråga .
Är det då verkligen en tillfällighet att det nästan alltid är samma staters flagga , som dessa fartyg seglar under ?
Varför finns det då ingen svart lista ?
Om osäkra och farliga flytande likkistor färdas i europeiska farvatten , varför säger man då inte , liksom i andra sammanhang , att dessa inte får komma in i europeiska farvatten och inte får anlöpa europeiska hamnar ?
Alltså skulle jag gärna i er åtgärdslista för sommaren också vilja ha en total granskning av alla tankfartyg , som för närvarande färdas i europeiska vatten , och jag skulle också gärna vilja veta det senaste läget i fråga om vad Europeiska unionens medlemsstater nu faktiskt har skrivit under och genomfört i fråga om IMO-bestämmelser ( Internationella sjöfartsorganisationen ) och konventioner , ty där finns det också alltid en fördröjning .
Det som skedde med Erika var inte något slarv , utan från min synpunkt sett en kollektiv , brottslig ansvarslöshet , och vi i parlamentet har under de närmaste månaderna möjlighet att med hjälp av en sak bevisa om vi menar allvar : Det är hamnarnas uppsamlingsanläggningar , där det handlar om medlemsstaterna .
Vi kommer då att ses och tala med varandra igen , och jag hoppas att vi då alla är av samma uppfattning som i dag !
Herr talman , fru kommissionär !
Jag anser att den beklagansvärda händelsen med Erika i själva verket , så som man har påpekat här i eftermiddag , bör bli en definitiv vändpunkt som markerar före och efter den här typen av olyckor i Europeiska unionen , där det sedan 1967 har inträffat sjutton olyckor med stora oljetankfartyg , det vill säga mer än en olycka vartannat år .
De sociala och ekonomiska skadorna , som vi redan har talat om här i dag , både vad gäller en försämrad sysselsättning och försämrade resurser inom fiske och turism , är av den omfattningen att de mer än väl motiverar ett beslutsamt och övertygande agerande från gemenskapsinstitutionernas sida .
Även jag , fru kommissionär , vill tacka för kommissionens snabba reaktion på denna händelse och de åtgärder man nu vidtar och de som är på gång .
Och jag litar på att dessa åtgärder inom de närmaste månaderna leder fram till ett tydligt och övertygande rättsligt instrument - eventuellt ett direktiv - som en gång för alla sätter stopp för dessa pirater på 2000-talet , som berövar oss alla på havets rikedom och skönhet .
Jag skulle vilja göra ett påpekande beträffande en av de åtgärder som kommer att vidtas och som har påtalats av kommissionären och av flera av mina kolleger .
Det gäller dubbelskrovet , som innebär att lasten inte har kontakt med ytterskrovet , det vill säga skrovsidan mot sjön .
Fru kommissionär , det finns många experter som anser att dubbelskrovet inte är tillräckligt säkert och i stället rekommenderar ett så kallat " ekologiskt skrov " , där havsvattnet vid en eventuell olycka tränger in i tankarna och gör att oljan , på grund av trycket , förs över till andra tankar .
Jag anser , fru kommissionär , att det är dags att vi röstar på de säkraste tekniska åtgärder som finns .
Därför anser jag att vi inte får nöja oss med att kopiera en lagstiftning som gäller i andra länder .
Jag anser att vi kan och bör förbättra den lagstiftning som finns på området .
Varje analys av kostnader och vinst där man beaktar de totala skadorna på människorna och miljön till följd av dessa olyckor , kommer att ge oss rätt .
Herr talman , fru kommissionär , kära kolleger !
Jag skulle först och främst önska att vi gläder oss över vårt förfarande .
Det gör det möjligt för oss att slutligen lägga fram en gemensam resolution - efter det att alla politiska grupper har samlat sig för att uttrycka vad alla känner .
Under dessa tragiska omständigheter tror jag att det vore en missuppfattning och en skam om vi talade med flera olika röster , principiellt sett .
Det faktum att parlamentet i dag lägger fram en resolution med en enda röst - vi kunde konstatera de föregående talarnas samsyn - tror jag utgör ett tillfälle för oss parlamentariker att sätta press på ett antal regeringar , som tvekar och ägnar sig åt undanmanövrar , och jag tror att det är en mycket stark politisk handling som vi lägger i kommissionens händer för att förbereda ett europeiskt maritimt område .
Jag tror att det står helt klart - och det är den första slutsatsen man kan dra av Erikas katastrof - att allmänheten inte skulle förstå varför man antar bestämmelser för choklad men inte för transporter till havs .
Allmänheten skulle inte förstå varför man talar om ett gemensamt rättsområde , att man talar om ett gemensamt luftområde , att man talar om ett gemensamt järnvägsområde och en gemensam marknad , men inte om ett maritimt område .
I dag tror jag att det är ett arbete som måste inledas med en bestämd vilja till resultat , konkreta resultat .
Kommissionären pekade på tre stora avsnitt som bör utvecklas : en modernisering av vår lagstiftning , så att vi kan ta fram normer .
Till min stora tillfredsställelse noterade jag för övrigt att t.o.m. de euroskeptiska grupperna , som förespråkar staternas suveränitet , vädjar till Europa att fastställa bestämmelser , och jag tror att EU är rätt nivå för det .
Ibland reglerar vi saker som i stor utsträckning skulle kunna regleras på en lägre nivå .
På det här området bör vi ge ett svar till allmänheten .
Det är mycket viktigt och alla måste känna sig berörda , för när allt kommer omkring är vi internationellt sett inte mer än en halvö .
Det krävs således uppföljningsregler .
Efter en modernisering av vår lagstiftning måste vi också inrätta systematiska kontroller och slutligen tillämpa principen om förorenarens / den betalningsskyldiges ansvar , vilket självklart är en förebyggande princip .
Jag skall strax avsluta , men jag vill också säga att jag har lämnat en förfrågan till utskottet för transport och turism om en offentlig utfrågning , för att vi direkt skall kunna följa upp ärendet Erika och förse framtida reflektionsarbeten med nytt underlag .
Jag hoppas att alla politiska grupper kommer att stödja vår förfrågan om en offentlig utfrågning .
Herr talman !
Oljetankern Erika , vars ägandeförhållanden döljs av brevlådeföretag på Malta och kanske Italien och Grekland , hyrd av TotalFina för transport av olja , förliste utanför den bretagniska kusten med alla katastrofala följder det medfört .
Konsekvenserna för miljön , den europeiska havsmiljöns flora och fauna är enorma .
Orsaken till katastrofen måste sökas i oljetankerns försvagade struktur .
Folk tvivlar således på säkerheten för fartyg som transporterar farlig eller förorenande last .
Den internationella maritima organisationen har utgivit en internationell reglering för detta .
Stater kan utföra hamninspektioner .
I Europa är lagstiftningen strängare och man måste , är förpliktigad , att kontrollera 25 procent av de inlöpande fartygen enligt direktivet port-state control .
Men det verkar som om inte en enda medlemsstat uppnår denna procentandel på grund av brist på inspektörer .
Det står helt klart att det inte råder brist på lagstiftning .
Jag tror att kommissionären har alldeles rätt i det .
Det som fattas är tillämpning av den redan befintliga lagstiftningen .
Men hur skall det nu gå till när vi faktiskt har brist på inspektörer , ärade Europeiska kommission ?
Kan kommissionen försäkra att direktiv 93 / 75 om minimikrav för fartyg som anlöper eller avgår från gemenskapens hamnar med farligt eller förorenande gods verkställs på ett korrekt sätt i alla medlemsstater ?
Borde inte kontrollen över verkställandet skärpas ?
Skulle det inte vara lämpligt att på kort sikt , enligt exemplet från Rotterdam , börja kontrollera enligt ett poängsystem , där till exempel fartygets ålder räknas in , om det är enkelväggigt eller dubbelväggigt , om det seglar under bekvämlighetsflagg .
Kort sagt , kontroll av äldre fartyg under internationell standard skall ha högre prioritet än fartyg som uppfyller alla kvalitetskrav .
Erika byggdes av ett japanskt skeppsvarv , enkelväggigt .
För närvarande finns ytterligare fyra systerfartyg i trafik .
Bygget stoppades då för tiden på grund av att faran för rostbildning var extra stor för den typen av fartyg .
Vissa av dem seglar också under maltesisk flagg .
Nu väntar vi på nästa olycka .
Borde det inte vidtas några sanktioner , som kommissionären sade , mot klassificeringssällskapet ?
RINA har för närvarande fått dåligt rykte .
Malta är på väg att inleda anslutningsförhandlingarna .
Jag anser att Europeiska unionen kan bevilja Malta inträde endast om det finns garantier för att den maltesiska flaggan i fortsättningen kommer att segla prickfritt .
Mina damer och herrar !
Jag skulle uppskatta om ni ville visa litet bättre disciplin , för vi börjar bli försenade , och denna försening kommer att gå ut över den tid som är avsatt till frågestunden med frågor till kommissionen .
Herr talman !
Strax innan jag gick ned i kammaren fick jag ett e-mail med en ganska känsloladdad beskrivning från en svensk kvinna som hade valt att tillbringa nyårsaftonen vid den franska kusten i Bretagne i stället för att vara hemma och fira med sina släktingar .
Liksom många andra hundratals frivilliga hade hon sett förstörelsen , tvättat fåglar och städat upp efter de ansvariga som inte fanns vid kusten de kvällar och nätter , när de verkligen skulle ha behövts där .
Som så många andra , undrar även jag var de ansvariga finns .
Var finns redarna och transportbeställarna när dessa katastrofer inträffar ?
Kanske vore det dags för oss att börja fundera över att inrätta en gemensam miljöbrottsmyndighet , som skulle kunna ta upp denna typ av brott .
Det är inte första gången vi ser oljeutsläpp , avsiktliga eller oavsiktliga .
( Talmannen avbröt talaren ) Jag skulle vilja tacka Grossetête och hennes kolleger för att de har lagt fram detta förslag för parlamentet .
Brittiska massmedia har rapporterat mycket om miljökatastrofen då Erika sjönk utanför Bretagne och läckte ut 10 000 ton olja .
Trots att Storbritannien och Frankrike har haft sina meningsskiljaktigheter på senaste tiden kan jag försäkra er att mitt land känner stort medlidande med alla de drabbade .
TV-bilderna av den skada er kustlinje och ert djurliv , särskilt fåglar och det redan tynande fiskbeståndet , har lidit fick oss att minnas liknande katastrofer i Storbritannien , såsom Torrey Canyon 1967 , och har fått många britter att ställa upp med frivilligt arbete .
Jag välkomnar dessa gemensamma ansträngningar att reparera skadan .
Det är tydligen ett problem för hela EU : s kustlinje som kommer att kräva fantasifulla lösningar .
I stället för att låta de mest drabbade områdena och försäkringsbolag som Lloyds i London bära kostnaderna för dessa katastrofer måste vi utveckla nya tekniker för att återvinna mycket mer än 10 procent av den förlorade oljan från havet .
Eftersom försäkringsmarknaden betalar räkningen för närvarande finns små ekonomiska incitament för detta .
I slutändan måste den som förorenar betala .
Dessutom måste vi bygga vidare på rådets direktiv om genomdrivande av internationella normer för fartygssäkerhet och förebyggande av föroreningar genom att säkerställa att målet att 25 procent av de fartyg som anlöper EU : s hamnar skall kontrolleras uppfylls och att kontrollerna håller hög standard .
Dessutom anser jag , även om jag inte är emot att fartygens ägare registrerar sina fartyg i vilket land de vill , att en striktare tillämpning av internationella bestämmelser fordras .
Snarare än att förbjuda bekvämlighetsflagg , vilket skulle vara ett brott mot varje suverän stats rätt att ha en handelsflotta , måste nationella sjöfartsmyndigheter i enlighet med 1995 års EG-direktiv om hamnkontroll pålägga utflaggningsländer som inte uppfyller sina åtaganden enligt internationella avtal effektivare sanktioner .
Jag hoppas verkligen att kommissionen och rådet , speciellt under det franska ordförandeskapet senare i år , kommer att titta noggrant på dessa alternativ och jag rekommenderar helhjärtat parlamentet att anta denna resolution .
Herr talman !
Det är nästan kusligt att i dag återigen stå här , med regelbundna mellanrum sedan nästan 10 år , på grund av en olycka som orsakats av människohand och brist på mänskligt förnuft , och inte på grund av force majeure .
Där ute väntar de drabbade .
De vill ha svar .
De vill inte ha några fler löften , som vi sedan ändå inte håller , de vill inte ha några ansträngningar , som vi sedan ändå inte slutför .
Befolkningen frågar med all rätt : Hör våra regioner nu till dem som slutgiltigt gått förlorade ?
Vem skall ge oss några nya arbetstillfällen ?
När skall upphovsmännen äntligen begripa att skonandet av resurserna inte är någon fritidssysselsättning , inte någon fråga för ett enda system eller för en ny arbetsgrupp , utan en gemensam europeisk utmaning ?
Därför , fru Palacio , är er handlingsplan mycket välkommen .
Lika väsentligt är följande : Det är viktigare att förebygga än att bota .
Men man måste också ha kunskaperna .
Insatserna som gjordes av det tyska allroundfartyget Neuwerk - det ligger just utanför min husdörr i Cuxhaven - innebar en snabb europeisk grannhjälp .
Ett uttryckligt tack gäller de svåra insatser som gjordes av allt manskap .
Man samlade värdefulla erfarenheter , men insåg också att vi enbart med hjälp av modernaste teknik inte kan bemästra sådana miljökatastrofer .
Vi kräver alltså med all rätt bättre kontroller , påföljder och säkerhetsåtgärder .
I snart tio år har jag här i parlamentet kämpat för en europeisk miljökustbevakning .
Frågan är lika aktuell som någonsin .
Jag kommer också i fortsättningen att ställa upp , och gemensamt med andra satsa på att åstadkomma förbättringar och logiska koncept inom ramen för ett europeiskt respektive internationellt samarbete .
( Applåder ) Herr talman !
Jag vill börja med att uppriktigt tacka för alla initiativ , inte bara från de olika grupperna , av Grossetête och av Europeiska folkpartiets grupp ( kristdemokrater ) och Europademokraterna , utan även från Wurtz och Gruppen Europeiska enade vänstern / Nordisk grön vänster , till denna debatt som har gjort att vi har kunnat föra en viktig diskussion i positiv anda .
Min avsikt är att lägga fram ett meddelande före utgången av mars månad , och det är möjligt att det kommer att innehålla lagtexter , det vill säga ändringar av konkreta direktiv så att en diskussion kan föras i rådet och i parlamentet .
Jag skulle vilja påstå att det här i själva verket inte bara handlar om ett miljöproblem ; det är ett omfattande miljöproblem , men det är också ett omfattande socialt problem ; det finns män och kvinnor som är beroende av fångst av fisk och skaldjur , av tjänstesektorn eller turistsektorn i dessa kustområden ; det är områden som är utsatta ur miljösynpunkt , men även utsatta vad beträffar den sociala utvecklingen och den territoriella jämnvikten .
Därför måste vi vara särskilt försiktiga så att vi i den mån det är möjligt undviker att en situation som denna uppstår igen .
Roth-Behrendt sade att ingenting har gjorts .
Jag tror nog att kommissionen tidigare har gjort en del , men ännu mer måste göras .
Beviset på detta är att nordamerikanerna , efter Exxon Valdez , inom ett år antog en lagstiftning som var extremt sträng och extremt hård , och som innebär en risk att man , som jag redan har påpekat , omdirigerar de båtar hit som inte accepteras av de nordamerikanska hamnarna .
I Europa har vi , sedan Amoko Cadiz eller Urquiola vid den spanska kusten år 1976 eller Torrey Canyon samma år , eller sedan alla andra fall som har förekommit , börjat lagstifta på allvar sedan år 1994 och 1995 , och i synnerhet på senare år .
De senaste åren har man dessutom poängterat säkerheten vid passagerartransporter .
Sådan är verkligheten .
Enligt min uppfattning måste vi nu göra viktiga och angelägna insatser för att bemöta de nya problemen , som även härrör sig från den nordamerikanska lagstiftningen , där man poängterar säkerheten vid transport av farligt gods inom sjöfartssektorn .
Mina damer och herrar , jag har tagit upp en rad frågor som vi kan gå in på mer i detalj , om ni vill , i samband med att jag infinner mig i det utskott som berörs av frågan , eller annars i samband med att jag lägger fram konkreta initiativ de närmaste månaderna .
Min avsikt är - och det är något jag vidhåller - att vi påbörjar diskussionen i slutet av mars , en tidpunkt som sammanfaller med ett ministerråd , och att vi , givetvis innan det portugisiska ordförandeskapets period är till ända , får ett diskussionsunderlag .
Bekvämlighetsflaggen är ett problem , men det är inte det enda .
Rumänien är inte ett land med bekvämlighetsflagg , men man har ändå en mycket hög felkvot vid inspektioner .
Ännu högre än länderna med bekvämlighetsflagg .
Malta och Cypern har begärt inträde i unionen .
Vi måste ställa höga krav i den här frågan och nu pågår förhandlingar om detta .
Det kommer att leda till att vi får ompröva Europeiska unionens register och ta upp det välkända problemet , som säkert kommer att dyka upp igen , vilket syftet är med ett gemenskapsregister .
Även om jag tror att det skulle vara svårt , bör man utföra en granskning av de register som finns i Europeiska unionens länder .
Vad beträffar kontrollerna , så är själva kärnfrågan , det vill säga det första man måste ta reda på , hur den lagstiftning som vi förfogar över har fungerat , precis som Hatzidakis påpekade .
Vi har ju redan en lagstiftning .
Enligt den information som kommissionens tjänsteenheter tillhandahållit mig har lagstiftningen i många medlemsstater inte tillämpats i tillräcklig utsträckning , på grund av brist på personal , resurser och inspektörer .
Problemet är inte att endast 25 procent kontrolleras , utan snarare hur urvalet går till , hur man hittar de fartyg som utgör den största risken , utifrån fartygens ålder eller utifrån flaggens tidigare riskfaktor .
Tyvärr gömmer sig dessa 25 procent bakom flagg som de vet kommer att uppfylla kraven : inspektionerna går då snabbare och arbetet är lättare att utföra .
Därför måste man , förutom att vidta förändringar , även vidta åtgärder för att undersöka vad som redan görs , förutom några tilläggskrav beträffande granskningarna , i synnerhet i förhållande till de olika fartygens ålder .
Där finns SOLAS ( Internationell konvention om säkerhet för människoliv till sjöss ) och MARPOL ( en internationell konvention om förhindrande av havsföroreningar från fartyg ) , två avtal inom ramen för Internationella sjöfartsinspektionen , som bör göras obligatoriska i unionens samtliga stater så att man sedan kan kontrollera hur de tillämpas .
Vad beträffar unionens inspektörer , anser jag att subsidaritetsprincipen motiverar att man godkänner att medlemsstaterna utför dessa inspektioner , vilket inte hindrar att kommissionen kontrollerar att staterna utför sin uppgift på rätt sätt .
Slutligen vill jag poängtera ansvarsfrågan .
Inte bara beträffande maxbeloppen som jag anser bör vara jämförbara med de nordamerikanska .
Vi har fastställt 180 miljoner dollar ; i Förenta staterna talar man om 1 000 miljoner dollar som ett tak för skadeersättning .
Jag anser att vi bör höja det aktuella beloppet , så att vi närmar oss de nivåer som finns i Förenta staterna , men att vi även bör kräva en omprövning av totalsumman för försäkringarna av fartygen , och därmed rederiernas ansvar , och låta ansvaret även omfatta dem som chartrar fartygen , ägarna av lasten .
Så länge man inte utkräver något ansvar av de som äger lasten , mina damer och herrar , så kommer dessa problem enligt mig inte att kunna lösas .
Det var allt , jag skall inte breda ut mig mer än såhär .
Vi kommer att få andra tillfällen att diskutera detta .
Men det är utan tvekan så att vi , som någon talare sade - och jag tackar för era inlägg som alla varit positiva och relevanta - måste förhindra att vi inom ett , två eller tre år åter står här och säger att vi inte har gjort det vi bör .
För min del kan jag , efter att ha diskuterat det med de övriga kommissionärerna , säga att kommissionen är beredd att inför parlamentet och rådet lägga fram de lagstiftningsåtgärder , ändringar och direktiv som krävs för att tillförsäkra oss den högsta möjliga säkerhetsnivån .
Detta förutsätter en politisk vilja från parlamentet- och jag ser att jag kan räkna med den - liksom även från ministerrådet .
Tack så mycket , fru kommissionär .
Vi har med glädje noterat er samarbetsvilja .
Jag har fått 8 resolutionsförslag i enlighet med punkt 2 i artikel 37 i arbetsordningen till följd av kommissionens uttalande .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum på torsdag kl .
12.00 .
 
Stormar i Europa Nästa punkt på föredragningslistan är kommissionens uttalande om stormarna i Europa .
Jag överlämnar ordet till Barnier som företrädare för kommissionen .
Herr talman , mina damer och herrar ledamöter !
Ni har just talat om de mänskliga , miljömässiga och sociala konsekvenserna av det oljebälte som än en gång har drabbat de franska kusterna .
Och vi kommer nu - vilket gläder mig personligen - att tala om konsekvenserna av en historisk storm , en verklig orkan som också och samtidigt drabbade Frankrike , men även Förbundsrepubliken Tyskland och Österrike .
Mina damer och herrar !
När man talar om konsekvenserna av olyckor och oväder av det här slaget , handlar det inte endast om skador på miljön och kulturarvet .
Då talar man också om , vilket även jag vill göra , vilka konsekvenser stormarna liksom oljebältet får för alla de kvinnor och män , vilket Loyola de Palacio sade för en stund sedan , alla de familjer som verkligen , det kan jag intyga , har blivit varaktigt chockade , skadade , märkta , missmodiga , och när det gäller de allra svagaste , förtvivlade .
Mitt intryck är att det här i dag uttrycks en europeisk solidaritet och att denna solidaritet tar sig uttryck i ord om moraliskt stöd , men att den framför allt är en mänsklig solidaritet .
Och jag vill uttrycka detsamma å hela kollegiets vägnar , och i synnerhet å de kollegers vägnar som varken glömmer var de kommer ifrån eller sitt medborgarskap ; Franz Fischler för Österrike , Michaela Schreyer och Günther Verheugen för Tyskland samt Pascal Lamy och jag själv för Frankrike .
Denna solidaritet åtföljer den som redan har markerats av dessa länders nationella myndigheter och av en fantastisk generositet och frivilliga insatser .
Och eftersom vi talar om Europa , vill jag också hylla spontaniteten och tjänstvilligheten hos frivilliga från offentliga företag som elleverantörer , telebolag , brandkårer och vägförvaltningar , som kom spontant från hela Europa för att hjälpa till att få igång trafiken igen , och på vissa håll elektriciteten och telefonnäten .
En del familjer i vissa franska regioner , mina damer och herrar , har inte kunnat ringa eller inte haft ström förrän för ett par dagar sedan .
På begäran från ordförande Romano Prodi har kommissionen haft ett första samtal om den här frågan i sin helhet , en diskussion under kommissionens första sammanträde för i år .
Och jag vill därför , vilket ordföranden har bett om , delge er resultatet av vårt arbete för att komma fram till vad unionen kan bidra med inom ramen för förordningarna och budgeten när det gäller återuppbyggnaden av det ekonomiska , sociala och kulturella arv som har skadats , efter att ha uttryckt vår mänskliga och moraliska solidaritet .
Mina damer och herrar !
Kommissionen kommer att uppbåda alla instrument som står till vårt förfogande för att hjälpa de berörda medlemsstaterna med återuppbyggnaden och ge stöd till drabbade personer eller företag , för att åtfölja och komplettera det stöd och den hjälp som nationella och regionala myndigheter redan har fattat beslut om .
Ni vet att kommissionen förfogar över flera instrument , flera redskap som kan ge bidrag till sanerings- och återuppbyggnadsinsatserna , och vi räknar med att utnyttja alla dessa instrument med en lika stor viljekraft som Loyola de Palacio uttryckte när hon talade om lärdomarna av Erika-katastrofen .
När det gäller strukturpolitiken , kommer jag personligen att granska hur vi kan utnyttja de beslut som nu fattas om den nya generationen ekonomiska utvecklingsstrategier - som kommer att tillämpas under de sju kommande åren , och hur de redan beviljade totalanslagen - särskilt för landsbygds- , industri- och tätortsregioner som genomgår en omställning och för fiskeområden , dvs. de regioner som omfattas av mål 2 - kan bidra till återuppbyggnaden .
Områdesindelningen för mål 2 har fastställts av kommissionen efter samråd med de olika regeringarna .
För Tyskland fattade kommissionen beslut i december , och just i dag har kommissionen fastställt mål 2-kartan , inte bara för Luxemburg och Sverige , utan också för Frankrike och Österrike .
För Frankrike , där skadorna objektivt sett är störst , finns det totalt 5,4 miljarder euro att tillgå i det nya mål 2 under perioden 2000-2006 .
En första analys som har gjorts av kommissionens enheter visar att 70 procent av de personer som har drabbats av ovädret kommer att få stöd från mål 2 , utifrån en finansiell fördelning i proportion till den befolkning som är stödberättigad .
De 69 olycksdrabbade franska departementen skulle därmed kunna få omkring 4,1 miljarder euro under de sju kommande åren .
För Tyskland och Österrike är de motsvarande totala beloppen 3 miljarder euro för Tyskland och 600 miljoner euro för Österrike .
Jag vill också erinra om , mina damer och herrar ledamöter , att de olycksdrabbade områden som inte finns med på den nya kartan - och tyvärr finns det också sådana - dvs. de som inte berörs av mål 2 , men som enligt den tidigare områdesindelningen var berättigade till mål 2 och mål 5b , också kommer att få tillgång till de anslag som finns tillgängliga för den nya programperioden , dvs. stöd under en övergångstid .
Jag vill således klart och tydligt påpeka att strukturanslagen i hög grad kan bidra till de olycksdrabbade områdenas ekonomiska sanering .
Det handlar givetvis inte om något katastrofstöd - ni vet för övrigt mycket väl att de blygsamma anslag som fanns tillgängliga i EU-budgeten för katastrofstöd avvecklades för två år sedan - det handlar i stället om ett återställande och en sanering på lång sikt , inom ramen för de program som är under förberedelse , och det är ur min synvinkel det viktigaste .
Programplaneringen för åtgärder och val av prioriteringar har , som ni vet , decentraliserats till varje enskild stat , och därför kommer varje regering att behöva fastställa sina prioriteringar och göra sina val utifrån de förutsättningar jag just nämnt .
Det blir troligtvis nya prioriteringar , med hänsyn till stormarnas eller oljebältets konsekvenser .
Det åligger de berörda ländernas regeringar att fördela gemenskapens finansiella stöd mellan de olika regioner som är berättigade till strukturstöd , och därmed att föreslå kommissionen de handlingsplaner som kommer att genomföras på plats .
Men för att ta ett exempel , för att vara mer konkret , vill jag erinra om att alla dessa program kommer att kunna finansiera de olycksdrabbade regionernas återställande av det historiska och kulturella arvet , deras ekonomiska aktivitetsområden , industri- och hantverksområden , det vägunderhåll som krävs för avsättning av råvaror och industriprodukter , infrastrukturen i hamnarna : handels- och fritidshamnarna ; de flygplatsinfrastrukturer som är viktiga för affärsresor och turism ; produktiva industriella investeringar ; stöd till företag ; det historiska och kulturella arvet av turistiskt intresse samt utbildning av behörig personal med stöd ur Europeiska socialfonden .
Kommissionen står således till medlemsstaternas förfogande , för att justera och på bästa sätt omstrukturera programplaneringen , och det gäller även , det vill jag understryka , dem som drabbades av andra oväder i början av december , i Danmark , Förenade kungariket och i Sverige .
Jag känner till att parlamentet antog en resolution den 16 december om den frågan .
Eftersom jag var där två gånger vill jag erinra om att detta också gäller Grekland , med anledning av konsekvenserna av jordbävningen i början av september och mål 1 i Sammanhållningsfonden .
Mina damer och herrar !
Min kollega Franz Fischler har samma strategi för landsbygdens utveckling .
Efter reformen av den gemensamma jordbrukspolitiken , som godkändes av parlamentet i fjol , kan åtgärder för landsbygdens utveckling för första gången samfinansieras av Europeiska utvecklings- och garantifonden för jordbruket ( EUGFJ ) , garantisektionen , i unionens alla landsbygdsområden .
Således kommer Frankrike att få 760 miljoner euro per år , Tyskland 700 miljoner euro och Österrike 423 miljoner euro .
Dessa stöd är tillgängliga för de olycksdrabbade regionerna , men utan den begränsade områdesindelning som jag är tvungen att tillämpa för mål 2 .
Bland de åtgärder som kan finansieras av EUGFJ , garantisektionen , vill jag nämna återställandet av den skadade jordbruks- och skogspotentialen , skogsåterväxten , infrastrukturerna på landsbygden , förebyggande och skyddande infrastrukturer , såsom hinder och varningssystem .
I det sammanhanget är skogsindustrins problem troligen det mest specifika , eftersom den blev särskilt drabbad av stormarna .
Vi kommer att ägna den en särskild uppmärksamhet , såväl ur ekonomisk som miljömässig synvinkel .
När det gäller virkeslagren vill jag säga att EUGFJ också kan stå för gemenskapens samfinansiering .
När det för övrigt gäller fisket , är det även möjligt att uppbåda strukturinstrumenten för samfinansieringar .
Frankrike har tillgång till 225 miljoner euro för perioden 2000-2006 .
Gemenskapens stöd kan bidra till att ersätta fiskare och fartygsägare för tillfälliga avbrott i deras verksamhet i händelse av oförutsedda händelser , och det under högst två månader per år .
Stöd från det finansiella instrumentet för utveckling av fisket ( IFOP ) är också tänkbart , möjligt att utnyttja för klassiska investeringsprojekt .
Jag tänker på vattenbruksanläggningar , kollektiva anläggningar , omstrukturering , fysisk planering av vattenbruk , utrustning för fiskehamnar , modernisering av fartyg .
Jag har redan förhört mig om de frågorna tillsammans med Franz Fischler .
Kommissionen vill slutligen betona att de statliga stöd som är avsedda att reparera de skador förorsakade av naturkatastrofer eller andra extrema händelser kan komma att anses förenliga med den gemensamma marknaden , givetvis efter samråd med min kollega Mario Montis enheter , och skulle då godkännas av kommissionen .
Redan nu kan således olika åtgärder sättas in , i fråga om energi kan det till exempel ske inom ramen för programmet för transeuropeiska nät för energi .
När det gäller transport av energi är jag väl medveten om att det finns många tekniska problem , i synnerhet transport av energi via högspänningsledningar .
Men eftersom jag minns den inte alltför avlägsna period då jag var miljöminister i Frankrike , när jag stred för en nedgrävning av ledningar , vill jag erinra om det som vissa av er sade för en stund sedan , nämligen att det är mycket billigare att förebygga än att rätta till i efterhand , på detta område liksom så många andra .
Jag skulle därför önska att medlemsstaterna när det är tekniskt möjligt främjar en nedgrävning av telegrafi- , telefoni- och elledningar , och att vi uppmuntrar dem till det .
Mina damer och herrar ledamöter !
Så långt presentationen av de gemenskapsinstrument som erbjuder ett stort antal mycket konkreta interventionsmöjligheter .
Europeiska unionen gör inte allt , och kommer inte att göra allt .
Men den kan göra mycket , under förutsättning att vi har förmågan att uppbåda dessa instrument , att ni informerar om detta och att medlemsstaterna kan fastställa sina prioriteringar och fatta sina beslut till följd av stormarna .
Det är således mycket viktigt att kammaren , liksom kommissionen , vidarebefordrar denna information och detta konkreta solidariska budskap till alla berörda parter samt berörda och drabbade människor .
Vad mig beträffar åtar jag mig att göra detsamma redan denna vecka , eftersom jag i övermorgon beger mig till två franska departement som blev hårt åtgångna av stormarna : la Charente-Maritime , drabbat av såväl orkanen som oljebältet , och la Creuse .
Jag kommer också att presentera dagens beslut om mål 2 .
I morgon , den 19 januari , kommer min kollega Michaela Schreyer att besöka en av de värst drabbade regionerna i Tyskland , Svarta Skogen i Baden-Württemberg .
Jag vill avsluta denna framställning genom att tacka för er förståelse , herr talman , och genom att ta upp ett ämne som ligger mig varmt om hjärtat och som är en av de lärdomar vi bör dra av dessa katastrofer , inte alltid , men ofta naturkatastrofer .
Vi är övertygade om att den här typen av katastrofer förstärker behovet av en bättre samordning inom unionen av de medel som finns i varje stat för gottgörelse , katastrofstöd och civilt skydd .
Kommissionen har redan en samordningsenhet på området för civilt skydd , vilken är placerad under min kollega Margot Wallströms ansvar .
Denna enhet har för övrigt fungerat väl när det har handlat om att hantera oljebältet , att hitta båtar , upprätta strandskydd och ta fram maskiner för att inom gränsen för det möjliga rengöra oljeindränkta fåglar .
Här har man uppbringat medel från elva europeiska länder , något man inte alltid känner till och något som motiverar den hyllning jag ville ge denna spontana solidaritet , som alla europeiska länder har visat .
Emellertid anser jag att vi måste gå längre än så .
Ordförande Prodi , Margot Wallström och jag själv är övertygade om att det krävs att man på ett mycket mer systematiskt sätt utvecklar en europeisk interventionsstyrka som stöds på befintliga nationella bestämmelser och på specialiserade enheter .
Dessa skulle kunna utgöras av brandmän , vaccinations- och civilskyddsenheter , spårhundar vid lavinolyckor och mycket mer och medlemmarna av en sådan styrka skulle vara kvar i sina respektive länder men följa en gemensam utbildning och träning , och de skulle vid behov kunna mobiliseras på Europeiska unionens territorium , till exempel som man såg i samband med stormarna och jordbävningen i Grekland , och även utanför unionen , som i Turkiet , Sydamerika och Centralamerika , till följd av de tragiska händelser vi alla känner till .
Det verkliga frågan är huruvida det är möjligt att upprätta en verklig europeisk civil skyddsstyrka .
Dit har vi ännu långt kvar i dag , även om Europeiska rådet i Helsingfors tog ett steg framåt i den riktningen och Margot Wallströms enheter arbetar på en utvidgad roll för " interventions- och spaningsstyrkan " .
För stunden har kommissionen självklart varken de mänskliga resurser eller ekonomiska medel som krävs för att kunna åta sig ett sådant uppdrag , men tillsammans med Margot Wallström och under Romano Prodis ledning anser vi att detta är en av de lärdomar som bör dras efter den senaste raden av olyckor - naturkatastrofer eller ej - med så tragiska konsekvenser .
Det skulle också vara , i fråga om effektivitet och politisk tydlighet , en symbol för vår föreställning om Europeiska unionen .
Vad mig beträffar har jag för avsikt att inom kollegiet framföra denna idé som en av de lärdomar vi bör dra av de senaste katastroferna .
Herr talman !
Under 1999 års sista dagar svepte oerhört våldsamma stormar fram , i huvudsak drabbades Frankrike , men också Tyskland , Spanien , Förenade kungariket och Schweiz .
Man har tyvärr kommit fram till 100 döda , varav 88 i Frankrike .
De mänskliga skadorna är enorma , men också den materiella förstörelsen ; offentliga anläggningar och privata egendomar har förstörts eller skadats allvarligt .
Miljontals hushåll har stått utan elektricitet , telefon och rinnande vatten .
Ekonomisk verksamhet har stått stilla .
Enbart i Frankrike uppskattar försäkringsbolagen redan nu kostnaderna för skadorna till 35 till 40 miljarder franc , dvs .
5 till 6 miljarder euro .
Denna naturkatastrof , som saknar tidigare motstycke , har mobiliserat alla tillgängliga krafter och framkallat solidaritetsyttringar både inom och utanför gemenskapens gränser .
Därför skulle jag här vilja tacka alla dem som kom för att ge en hjälpande hand till räddningstjänsterna och de offentliga myndigheter och företag som översvämmades av den omfattande uppgiften .
Till alla er : ett tack ur hjärtat för denna värdefulla hjälp .
När chocken väl har lagt sig och våra samhällens vitala funktioner har återupprättats , funderar jag , och jag uppmanar också kommissionen och rådet därtill , över möjligheten att inrätta en post för katastrofstöd i gemenskapens budget , för att vi skall kunna hantera den här typen av händelser .
De risker som hänger samman med väderkatastrofer får inte försummas , och inför konsekvenserna av sådana katastrofer och de snabba interventioner som då krävs , tror jag det vore bra om gemenskapen på nytt försåg sig med sådana medel .
Detta katastrofstöd , som en gång tidigare existerade , borde kunna undantas från de strikta regler som tillämpas för strukturfonderna .
Jag instämmer också i kommissionär Barniers förslag att successivt inrätta en europeisk civil säkerhetsstyrka - en idé han lanserade redan för några månader sedan - och som vi talade om , herr kommissionär , när jordbävningarna inträffade .
På min fråga om möjligheten att återupprätta gemenskapens katastrofstöd , måste svaret självklart bli ja .
Jag skulle sedan vilja ta upp de oändliga problem som uppstår för en sektor som är synnerligen drabbad av stormarna .
Det gäller skogsbruket , vars verksamhet i allra högsta grad har äventyrats av de skövlingar som ovädret orsakade i skogarna .
Man måste förstå att skogen inte endast har en landskaps- och miljödimension .
De utgör också en viktig socioekonomisk sektor i vissa regioner , som inte får försummas .
I Frankrike har mer än 120 miljoner kubikmeter träd rivits upp av vindarna .
Det utgör ungefär tre års full skörd för producenterna .
Konsekvenserna är omedelbara .
Vissa skogsbrukare har förlorat allt .
Hela skogspartier har skövlats , vilket inom några veckor kommer att skapa säkerhetsproblem och fordra en bekämpning av bränder .
Priserna har redan rasat till följd av den enorma tillgången på trä , på grund av den övermättade marknaden .
Infrastrukturerna kommer att utsättas för en osedvanligt tät ström av långtradare och transport- och truckfordon .
Under dessa omständigheter är det brådskande att återupprätta tillträdet till skogspartierna , att återställa markerna och utnyttja tekniska lösningar för att iordningställa lagerutrymmen , hålla uppe priserna på trä , och på längre sikt bör man med alla tillgängliga medel underlätta skogsåterväxten .
Detta är en rad åtgärder som det finns anledning att vidta , herr talman , och jag gläder mig åt kommissionärens påpekanden , i vetskap om att mål 2 inte kan erbjuda stöd till allt .
Médoc är till exempel inte berättigad till detta stöd , herr kommissionär , och därför önskar jag att EUGFJ kan ersätta mål 2 i det fallet .
Herr talman , herr kommissionär , mina kära kolleger !
De osedvanligt våldsamma stormarna som har rasat i flera olika europeiska regioner bör parlamentet inte betrakta som ett dramatiskt , fast tillfälligt och exceptionellt fenomen .
Stormarna och konsekvenserna av dem är faktiskt en politisk händelse av stor vikt .
Varför ?
Varför skulle det inte vara en exceptionell händelse ?
Först och främst för att man i dag vet att liknande klimatfenomen aldrig är helt oförutsägbara .
Man vet nu att den här typen av oväder ofta hänger samman med klimatförändringar och växthuseffekten , och det är frågor för vilka medborgarna förväntar sig att Europeiska unionen skall utveckla en övergripande strategi för studier och prognoser .
Men vad som också står på spel i det här fallet - och som är skälet till att detta är ett utomordentligt viktigt politiskt fenomen för oss - är Europas förmåga att vara det man ger sig ut för att vara : ett Europa nära medborgarna .
I dag innebär det givetvis att vi måste sända ett starkt solidariskt budskap till alla dem som drabbats av stormarna , de familjer som förlorat en nära anhörig - jag vill erinra om att vi beklagar att minst 90 personer har dött till följd av ovädret - till de hantverkare som har förlorat sina arbetsredskap , de jordbrukare som på några ögonblick förlorade år av arbete , och till alla dem som firade övergången till det 21 : a århundradet i kyla och stearinljusens sken .
I det avseendet gläder jag mig åt det arbete som de politiska grupperna har ägnat sig åt de senaste dagarna , för att nå fram till en gemensam resolution som jag hoppas kommer att antas i morgon .
Men på ett konkret plan , och bortsett från alla ord , måste denna solidaritet självklart ta sig uttryck i en stor finansiell kraftsamling , som gör det möjligt att återuppbygga skadade produktionsled och förstörda kommunikationsnät , och att helt enkelt åter ge befolkningen värdiga levnadsvillkor .
Jag har förstått att en del av de olycksdrabbade områdena är berättigade till gemenskapens strukturstöd , och att man kommer att göra allt för att uppbåda dessa medel så snart som möjligt .
Men tillåt mig säga att detta inte är tillräckligt .
Det är inte tillräckligt eftersom dessa oförändrade totalanslag riktas om till reparation av skador , vilket följaktligen bestraffar investerings- och utvecklingsprojekt som var planerade på lång sikt .
Och lösningen förefaller framför allt oacceptabel med tanke på vilket europeiskt politiskt ansvar vi har gentemot allmänheten .
Medborgarna skulle inte förstå varför Europeiska unionen kan frigöra omfattande stöd vid enstaka katastrofer för att hjälpa offren för naturkatastrofer i tredje världen , även om ett sådant stöd är helt och hållet välgrundat .
Om vi vill se till att medborgarna inte uppfattar Europa som en maskin som producerar krångliga och petnoga bestämmelser , måste vi ändra på allt detta .
Vi måste fundera över ett nytt finansiellt arrangemang , som gör det möjligt att i brådskande fall uppbringa tillräckliga medel .
Och mot bakgrund av den stora mobilisering av transporter och mänskliga resurser som vi fick se när tekniker kom från hela Europa , bör vi främja inrättandet av en europeisk civil säkerhetsstyrka .
Det är i olyckan som man får reda på vem som står en nära och som man värderar deras solidaritet .
Jag tror att man bygger upp medborgarnas Europa till det priset .
( Applåder ) Herr kommissionär !
Jag vill tacka för era uttalanden , särskilt de konkreta förslagen angående de olycksdrabbade som väntar sig oerhört mycket av Europeiska unionen , och av det stöd som vi kan ge dem .
Några dagar efter de hemska stormarna sände jag personligen en skrivelse till er , för att be er att försöka få den franska regeringen att justera mål 2-områdena , så att alla drabbade områden kan få mål 2-stöd , såväl i Frankrike som i andra länder .
Jag antar att det är gjort , eftersom ni inte talade om det .
Vi vet att man har alla svårigheter i världen att få stöd om man inte ingår i ett mål 2-område .
Det är således bättre att genast lösa det här problemet .
Ni vet också att det inte endast är ett kortsiktigt problem , utan även ett problem på medellång och lång sikt .
Jag skall förklara mig .
Jag var i Lorraine när de förfärliga stormarna skövlade omkring 20 procent av lövskogarna .
För vissa s.k. skogskommuner är skador på 20 procent en enorm förlust .
Vi vet till exempel att det krävs mellan 150 och 200 år innan ett träd uppnår mogen ålder .
Den förlust som drabbar dessa kommuner sträcker sig således inte endast över ett , två eller fem år , utan en mycket längre period .
De berörda kommunerna uppskattar att det rör sig om 40 år .
Jag anser följaktligen att det kommer att bli mycket svårt att med hjälp av bidrag kompensera dessa landsbygdskommuners intäktsförluster .
Den aspekten tror jag att vi måste bära med oss och inte glömma den när vi vidtar olika politiska åtgärder .
Det stämmer att skogssektorns problem är oerhört sammansatt .
Ni talade om att frigöra medel för virkeslagren , eftersom priset inte får sjunka .
Å andra sidan kommer även de kommuner som inte berördes av stormarna att lida skada , eftersom Office national des forêts ( ung .
Skogsvårdsmyndigheten ) har beslutat att frysa skogsavverkningen under fyra års tid .
De kommuner som inte har lidit förluster kommer således ändå att få se sina inkomster minska .
Detta säger jag för att visa er att problemet är ytterst invecklat , och jag vill än en gång tacka kommissionen för att den analyserar situationen så grundligt som möjligt .
Jag skulle också vilja uppmärksamma er på det faktum att det visserligen har inträffat en ekonomisk katastrof , men att de verkliga miljökatastroferna ännu inte har inträffat .
Det sade ni själv , herr kommissionär - stormarna är inte alltid naturkatastrofer , och vår bedömning är att de är ett första tecken på klimatförändringar .
Vi bör därför se över vår politik för att integrera denna omständighet .
Herr talman , herr kommissionär !
Frankrike befinner sig fortfarande i ett chocktillstånd efter den förfärliga katastrof som orsakade ett tiotal personers död .
Ingen sektor besparades : alla infrastrukturer ; vägar , luftfart , järnvägar , hamnar , el- och telefonnät ; bostadsområden , skolbyggnader , historiska monument , och ej att förglömma jordbruket och skogarna , som i många regioner har ödelagts .
Folk är som mest chockade där skadorna var störst , men ingen har gett upp inför detta olycksöde .
Redan de första dagarna , och än i dag , visas en enorm solidaritet och generositet .
Förtroendevalda , kommunalanställda , medborgare i Frankrike och hela Europa har mobiliserat sig för att hjälpa till .
Jag vill särskilt hedra de offentliganställdas engagemang och uppoffring - de har gjort generösa insatser med ett enda mål för ögonen : att hjälpa olycksdrabbade människor och återupprätta normala levnadsvillkor , elektricitet , transporter , telefon , utrustningar .
Genom att bevisa sin effektivitet i dessa prövande stunder , gjorde den offentliga sektorn sig gällande som en oundgänglig del av vårt samhällsliv .
Jag tycker att det uppmanar oss att reflektera , framför allt för att sätta stopp för den pågående avreglerings- och privatiseringsprocessen .
Det är självklart också brådskande att fortsätta att plåstra om sår , att förbereda återuppbyggnaden och restaureringen , och samtidigt ta lärdom av denna exceptionella katastrof .
Jag har lyssnat till Barnier och uppskattar hans förslag , men personligen ser jag ingen motsats mellan omedelbara och långsiktiga åtgärder .
Det verkar tvärtom som om situationen gör att förslaget från min grupp blir relevant nu i efterhand , dvs. förslaget att återupprätta en specifik budgetpost för naturkatastrofer inom unionen .
Det finns självklart också anledning att utöka strukturfonderna till förmån för de drabbade regionernas återuppbyggnad , bl.a. de medel som anslås till landsbygdens utveckling , livsmedelsåtgärder och skogsbruket .
Jag har särskilt noterat förslagen rörande mål 2 .
Man har framfört hypotesen att den här typen av katastrofer hänger samman med klimatförändringar , som uppstått till följd av människans aktiviteter i miljön .
Om detta bekräftas vore det också bra om unionen gör mycket större insatser för att få länderna att respektera åtagandena från Kyotokonferensen och prioritera planetens fortlevnad i stället för den ohämmade jakten på lönsamhet .
Herr talman !
Alla de som kom hit med bil , tåg eller flyg , har kunnat konstatera vidden av de skador som framför allt drabbat Frankrike till följd av orkanen , en orkan av en aldrig tidigare skådad styrka , som slog till mot Europa i slutet av förra månaden .
Vad kan Europaparlamentets ledamöter göra inför en katastrof av den omfattningen ?
Först och främst vill jag hedra alla mina kolleger , borgmästare och förtroendevalda , som varje dag har fått lugna människor , organisera solidaritetsarbetet och samarbeta med de offentliga tjänsteföretagen .
De har gjort sig väl förtjänta av sina medborgares förtroende .
Jag vill också tacka medlemsstaternas räddningstjänster och väpnade styrkor , som inom ramen för ett exemplariskt mellanstatligt samarbete kom för att stödja sina franska kollegers ansträngningar .
Jag skulle också vilja fundera över den paradoxala situation vi befinner oss i när det gäller katastrofstöd .
Hade denna katastrof ägt rum i Guatemala eller Turkiet hade vi genast kunnat ta gemenskapens budget i anspråk för att hjälpa offren , men i våra länder är inget sådant möjligt eftersom det saknas lämpliga budgetposter .
Vi måste också be kommissionen att inte hindra lokala myndigheter och staterna från att bistå de företag som har drabbats av katastrofen , dvs. att inte tillämpa gemenskapens konkurrensregler på ett alltför strikt sätt .
Jag tänker särskilt på de hårt drabbade fiskarna och mussel- och ostronodlarna .
Som ni sade herr kommissionär , måste de få ersättning för det påtvingade verksamhetsavbrottet , och de investeringar som måste byggas upp på nytt skall kunna få stöd genom det finansiella instrumentet för utveckling av fisket ( IFOP ) .
Vidare tror jag inte att en automatisk tillämpning av de fleråriga utvecklingsprogrammen ( FUF ) är på sin plats i olycksdrabbade kustområden .
Jag uppmanar därför kommissionen att avstå från det , för att i stället hjälpa dem som får sin försörjning av havet att göra de investeringar som nu är nödvändiga .
Herr talman , kära kolleger !
De stormar som härjade i Frankrike natten mellan den 26 och 27 december har som tidigare nämnts orsakat 90 döda och åsamkat skador för 75 miljarder franc , dvs .
11 miljarder euro .
Knappt tre veckor efter olyckan var tusentals människor fortfarande utan elektricitet och telefon , 500 000 hektar skogsområden och 100 miljoner kubikmeter träd hade förstörts och det historiska arvet hade också skadats , vilket det sorgliga exemplet Versailles slottspark vittnar om .
Inför en sådan katastrof förefaller det därför naturligt att den nationella och europeiska solidariteten kommer de olycksdrabbade och de mest berörda personerna till del .
Men i likhet med vad föregående talare har sagt , och vad ni , herr kommissionär , svarade min kollega Jean-Claude Martinez angående en annan tragedi - nämligen översvämningarna i sydvästra Frankrike i november månad - är det visserligen så att ni ser med oro på katastroferna , men det enda ni gör är att erinra om att budgetposten för hjälp vid naturkatastrofer har avvecklats .
Detta leder oss fram till en chockerande paradox , som framhölls av föregående talare , nämligen att det är lättare , mycket lättare , att hjälpa offren för naturkatastrofer utanför unionen än på unionens territorium .
Herr kommissionär !
Ni begränsar er till , och vi förstår er , att erbjuda oss den hypotetiska och avlägsna möjligheten att få strukturstöd enligt det nya mål 2 eller övergångssystemet för mål 2 och mål 5b .
Det var de ordalag ni använde i det skriftliga svaret till min kollega den 11 januari 2000 .
Jag har en kopia till ert förfogande .
Vi förstod mycket väl att ni inte kunde säga annat - inför den oansvariga attityd som inte endast är kommissionens utan också parlamentets - och att ni ingenting kan göra i brist på rättsliga och finansiella grunder .
Men för guds skull , jag ber er , och det säger jag utan någon som helst ilska gentemot er , presentera inte redan tidigare planerade stöd som hjälp till stormarnas offer , de är ju stöd som går inom ramen för en regionalpolitik som inte har någonting med detta att göra .
Inom ramen för en tilläggsbudget krävs det således att vi snarast återupprättar den budgetpost vi tilldelades för naturkatastrofer .
Vi måste utnyttja stödmedlen från toppmötet i Berlin , och vi måste ändra på den skogspolitik som bedrivs i de flesta av unionens länder , men det är ett annat problem .
Herr talman , herr kommissionär , mina kära kolleger !
Europa har vid detta millennieskifte utsatts för en hård prövning .
Först av allt vill jag uttrycka min djupa sympati med de familjer som försänkts i sorg av de oväder som härjade i Europa i december .
Stormarna är en miljökatastrof utan tidigare motsvarigheter för våra skogar .
Tillåt mig sända en särskild tanke till skogarna i min region , Lorraine , där skadorna var avsevärda .
Och jag vill gratulera de regionala myndigheterna , alla frivilliga och de offentliga företagen till deras exemplariska mobilisering .
Men tyvärr har de ännu inte sett ljuset i slutet av tunneln .
Det är Europas skyldighet att stödja dem och på så sätt komplettera de berörda medlemsregeringarnas insatser .
Jag välkomnar med nöje Barniers uttalande , liksom de åtgärder som kommissionen har aviserat .
Jag skall inte förbigå den ekonomiska dimensionen av frågan ; skogssektorn är ödelagd och en hel befolkning lider av de tragiska konsekvenserna .
Gemenskapens åtgärdsprogram för civilt skydd , vilket inrättades genom rådets beslut av den 9 december förra året , inleddes den 1 januari 2000 .
Jag vill be staterna att gripa tag i det tillfället : detta program måste fungera fullt ut .
Det har varit effektivt på vissa områden - och jag betvivlar inte att kommissionär Barniers uttalanden är ärliga - men jag beklagar att programmen för skogsbruket fortfarande ligger i sin linda .
I väntan på att medel frigörs på gemenskapsnivå , bör man prioritera ett materiellt stöd inom ramen för medlemsstaternas partnerskap .
Det är således brådskande att stärka skogssektorn och upprusta det så fort som möjligt .
Lån av skogsutrustning och tillhandahållande av behörig personal ingår också i ett sådant arrangemang .
En kommande utmaning blir att undvika växtskyddsproblem som hänger samman med att stora mängder trä överges i skogen , och att grundvattnet förorenas till följd av att det skapas lika betydande virkeslager .
Till sist är det absolut nödvändigt att bromsa utnyttjandet av avverkningsklara träd , och i stället främja köp av stormfällda träd .
Denna virkesförsäljning bör understödjas av en omfattande medial bevakning på medlemsstatsnivå .
Biståndet till uppsamling av trä utgör självklart bara ett första steg när det gäller att stödja återställandet av skogarna och den fysiska planeringen för landsbygden .
Jag uppmanar kommissionen att integrera detta i ett reflektionsarbete om förvaltningen av problemen efter katastrofen .
Det här är således ett sorgligt tillfälle för Europa att gripa tag i , så att dess skogrikedomar förnyas och skogarna därmed kan uppfylla sin uppgift att bevara vilda djur och växter och naturliga livsmiljöer samt sin roll i våra länders ekonomi .
För stunden krävs det således en solidaritet och ett samarbete mellan medlemsstaterna inför en ekonomisk och miljömässig katastrof .
Det är Europas sak att föreslå prioriterade åtgärder för att rädda skogssektorn , så att denna solidaritet verkligen blir meningsfull .
Orkanen " Lothar " måste ge oss anledning att överge vår princip att uteslutande återställa det som skadats , vilket också här diskuteras i främsta hand , och i stället tillämpa försiktighetsprincipen , där även de eventuella upphovsmännen skall ställas till ansvar .
De aktuella programmen måste påskyndas .
Åtagandet från Kyoto kan exempelvis inte genomföras med kommissionens nuvarande koncept .
Handeln med utsläppsrätter är enligt min åsikt omoralisk och löser inte problemet , utan skjuter bara upp det .
Hela skattesystemet måste på medellång sikt göras ekologiskt .
Genomförandet av uppgifterna i vitboken som rör förnybara energikällor , som skulle föra med sig en massiv minskning av växthusgaserna , måste påskyndas .
Allt som den nya kommissionen hittills har lagt fram i denna riktning , är inte på långt när tillräckligt , utan alltför litet !
Herr kommissionär , herr talman , mina damer och herrar !
Hittills har Lothar varit ett helt vanligt namn .
Men tyvärr har Lothar erhållit en beklaglig ryktbarhet .
Orkanen med samma namn svepte fram över Europa och krävde , framför allt i Frankrike och i Tyskland , men också i Schweiz , talrika offer , och efterlämnade en rågata med förödelse .
Vinden besegrade elmaster , tak , vägmärken och till slut också skogen .
Det rör sig ju bara om uppskattningar när vi nu hör att på kort tid ca .
120 miljoner fastkubikmeter träd fällts av stormen .
Jag har lyssnat mycket uppmärksamt på er , herr kommissionär , och jag välkomnar det också utomordentligt att ni kommer att ta en titt på katastrofen lokalt i Frankrike och Tyskland .
Om Schreyer nu under de kommande dagarna är i Schwarzwald , kommer den enskilde jordbrukaren eventuellt att fråga hur kommissionen nu skall kunna hjälpa honom .
Hur skall Europa kunna hjälpa mig ?
Vad säger ni då till skogsägaren , när hans skog eventuellt inte ligger i mål-2-området , om hans skog inte ligger inom 5b-området ?
Hur svarar kommissionen vid besöket på plats , när ni säger till skogsägaren att vi stöder vägbyggnad och dammar , vi vill bygga upp det kulturella arvet igen , vi vill komma med erbjudanden till turisterna etc ?
Att detta är välmenta råd .
Men jag kommer själv från en skogsfastighet i norra Tyskland , och jag kan tala om att vi i vår region redan nu märker dessa enorma skador .
Man fortsätter inte med den nödvändiga gallringen av skogen , skogarna sköts inte tillräckligt .
Vad vi ur kommissionens synpunkt absolut behöver , är också ett ja till de nationella stöden , så att vi inte senare åter talar om några konkurrenssituationer .
Herr talman , herr kommissionär , kära kolleger !
Tillåt mig att till att börja med visa på två fakta .
För det första : I början av 1999 jämnade Nato i frihetens namn Kosovo med marken med hjälp av bomber , med deltagande av de flesta medlemsstaterna i Europeiska unionen .
Nu försöker vi med gigantiska insatser åter få landet på fötter och hjälpa människorna där .
Detta med all rätt .
För det andra : I slutet av 1999 rasade oerhörda stormar och förde med sig död och förintelse över många landsändar inom EU .
Ropet på hjälp från de drabbade besvarades av kommissionen i Bryssel med en axelryckning .
Vi har inga medel och inga möjligheter , hette det .
Kära kolleger !
Detta är fel !
Ingen kan heller förstå det .
Och absolut inte den som känner sin existens hotad .
Människorna i Europeiska unionen förväntar sig solidaritet , även inom denna gemenskap .
Jag säger att de har rätt till solidaritet .
Europaparlamentet måste i nödens stund se till att de också får det .
Jag begär av kommissionen att den inte skall vara nödbedd utan gå offren för ovädret till mötes .
Kommissionen känner bättre till medel och vägar för hjälpen än alla lokala organisationer eller myndigheter .
Jag ber , kära kolleger , om ert stöd för att göra klart för kommissionen att det inte så mycket är möjligheterna att hjälpa som saknas , utan den goda viljan i många ämbetsrum i Bryssel !
Tillåt mig ytterligare ett påpekande : När det gäller stormens följder framgår detta mindre tydligt , men olyckan med tankfartyget utanför den franska kusten gör det helt klart att vi också i en annan fråga måste hjälpa kommissionen på traven .
Vi behöver inom Europeiska unionen snarast få regler beträffande miljöansvar .
Det går inte längre an att allmänheten får stå för de skador , som enskilda individer ofta orsakar med sina brottsliga förehavanden .
Vi måste göra upphovsmännen ansvariga för alla slags skador på vår miljö .
Då kommer exempelvis alla att överväga om de skall transportera olja i ett tankfartyg , som är på väg att brytas sönder .
När jag 1994 , för mer än fem år sedan , kom med i parlamentets utskottet för rättsliga frågor och den inre marknaden , fick jag ta över uppgiften som föredragande för området med miljöansvar .
Sedan dess väntar jag på ett initiativ från kommissionen , som också ger mig arbete .
Det är en skandal , som snabbt måste få ett slut , och jag hoppas att detta ärende inte skjuts upp än en gång i februari !
Herr talman , herr kommissionär !
Denna storm vid millennieskiftet bör få oss att tänka över problemen i grunden .
Det står klart att människan fortfarande inte är i stånd att undvika naturkatastrofer .
Det har alltid funnits och kommer alltid att finnas naturkatastrofer .
Naturligtvis behövs det solidaritet i detta sammanhang .
Det behövs säkerligen ett civilskydd över hela Europa , och det måste också inrättas en budgetpost för naturkatastrofer i EU : s budget .
Men - och det är det viktigaste - misstagen när det gäller förhållandet mellan natur och människa begås alltid av människan - även om de ofta görs över hundratals år - och aldrig av naturen , ty naturen kan inte göra några misstag .
Skadorna i detta sammanhang berodde på befolkningstätheten , på infrastrukturens utformning och i fråga om skogen naturligtvis också på de många monokulturerna .
Givetvis är jag positiv till att vi skall hjälpa så långt det är möjligt .
Men vid hjälpen skall man beakta att el- och telenät kanske i framtiden i större utsträckning bör läggas under jord .
Vi måste se till att vi får mindre kretslopp , och vid nyplanteringen av skog framför allt satsa på stabila blandskogar , och inte på monokulturer .
Den viktigaste diskussionen i detta sammanhang är emellertid klimatet .
Vi har hittills varit priviligierade i Europa , eftersom vi har Golfströmmen , och Golfströmmen fortfarande fungerar .
Amerika och Sydostasien har det mycket sämre ställt , vad gäller klimatet och stormarna .
Vi har lyckligtvis Golfströmmen .
Men vi lider liksom de andra också av växthuseffekten .
Den har - hur svårt det än är att demonstrera klimatförändringen med hjälp av räkneexempel - delvis åstadkommits av människorna .
Vi måste i större utsträckning iaktta direktiven från miljökonferensen i Kyoto .
Vi måste minska på koldioxidutsläppen , börja använda förnybara energikällor och i detta sammanhang generellt fråga oss , hur Europas skogar mår .
Herr talman !
Jag anser att det i första hand är offren vi bör beklaga .
Förlusterna är oersättliga .
För det andra välkomnar vi solidariteten de franska provinserna och medborgarna emellan , och övriga länders solidaritet med Frankrike som är det land som har drabbats hårdast .
Eftersom jag inte har så lång tid på mig , herr talman , vill jag endast ta upp två aspekter i vår resolution .
Den första tycker jag att kommissionären indirekt erkänner i sitt anförande , när han ställer sig frågan om det rör sig om naturkatastrofer eller ej .
Experterna blir ju ständigt mer övertygade om att det finns ett samband mellan klimatförändringarna och människornas agerande i allmänhet och det ökade antalet naturkatastrofer på senare år .
De senaste tio åren har temperaturen stigit mer än den hade gjort under den resterande delen av århundradet .
Därför bör Europa tydligt ta ställning för Kyotoprotokollet och komma med konkreta förslag .
Den andra aspekten är att det var jag som var föredragande för civilförsvaret i Europa , och jag är helt enig i kommissionärens förslag att upprätta en europeisk civilförsvarsmakt .
Dessutom bör man använda sig av en budgetpost utöver de vanliga , precis som en katastrofsituation är något utöver det vanliga .
Först av allt skulle vi vilja uttrycka vår medkänsla med alla de familjer och samhällen som har förlorat medlemmar i denna fruktansvärda tragedi .
Det är faktiskt förlusten av liv som gör denna speciella katastrof extraordinär med europeiska mått .
Det är beklagligt att vi inte har några verktyg för att ge bistånd i sådana här situationer .
Jag vill tacka kommissionären för hans innehållsrika uttalande i frågan och hans förslag att vi faktiskt skulle kunna organisera oss på europeisk nivå för att ge bistånd till medlemsstater och regioner som upplever liknande tragedier .
Detta är viktigt .
En andra sak vi bör komma ihåg är att vi hade en budgetpost tidigare .
Den var mycket liten .
Den räckte inte till mycket men den missbrukades flera gånger av ledamöter av denna kammare som föreslog åtgärder när katastroferna inte ens var stora .
Medlemsstaternas tjänstemän och ministrar kom till Bryssel , viskade med kommissionen , fick några euro och en politisk poäng genom att de hemförde stöd till sina valkretsar .
Så det var inte många som sörjde att denna budgetpost avskaffades .
Jag tror att vi bör återinföra denna budgetpost .
När vi hade jordbävningen i Grekland , som var en stor katastrof , hade inte gemenskapen något instrument för att visa grekerna sitt medlidande och sin solidaritet .
Detsamma gällde när översvämningarna drabbade Frankrike , och detsamma händer nu igen .
Dessa katastrofer är stora , vi borde ha ett instrument men vi har det inte .
Vi bör återinföra detta instrument och göra reglerna strikta , så att vi bara använder detta speciella instrument i situationer då allvarliga katastrofer inträffar .
Vi kan spara det från år till år och tillse att vi har ett instrument för att handskas med stora olyckor när de inträffar .
I Irland var det inte så illa den här gången , även om vi har haft många allvarliga stormar på Atlanten .
Vi hade översvämningar i Irland också och jag vill ge uttryck för min medkänsla med de människor i Irland som drabbades av dessa .
Mina kära kolleger !
Det får inte bli så att var och varannan bland oss tappar minnet .
Det stämmer att kommissionen och parlamentet fattade ett gemensamt beslut , vilket syftade till att avskaffa budgetposterna för katastrofhjälp .
Det stämmer att det finns mycket europeiska pengar - kommissionär Barnier har pekat på att han kommer att utnyttja artikel 30 i arbetsordningen om landsbygdens utveckling för ostronodlingarna och jordbruket ; artikel 33 för skogsbruket ; undantagen till konkurrensreglerna i artikel 87.2 i fördraget för företagens del samt strukturfonderna för offentliga anläggningar .
Ändå kvarstår det faktum att det i dag inte uppbringas ett enda öre mer än vad som skulle ha tilldelats före stormen , för att uttrycka en konkret och aktiv solidaritet .
För staterna gäller det helt enkelt att agera kommunicerande kärl och ta från ett ställe för att ge till någonting annat .
Detta är otillräckligt , och därför gläder det mig personligen att Barnier tog upp den idé som ligger mig varmt om hjärtat , en idé jag för övrigt framförde när jag uttryckte mina önskningar till pressen i Bordeaux , nämligen inrättandet av en förstärkt politik för ett europeiskt civilskydd .
Jag tror att medborgarna måste uppleva våra omedelbara åtgärder som påtagliga , om vi vill att det för oss så eftersträvansvärda europeiska medborgarskapet skall existera , och om vi vill att det mandat som vår talman Fontaine har ställt upp skall bli verklighet , dvs. att unionen och Europas medborgare skall närma sig varandra .
Jag tror därför att en europeisk civil säkerhetsstyrka borde vara något för oss att sträva efter ; att vi upprättar en formering av blå baskrar för civil säkerhet som skall vara närvarande på platser med svårigheter - inom unionen för att vi i dag inte har någon katastrofstrategi , men vid behov också utanför unionen , till exempel i Venezuela eller andra länder .
Jag vill också säga kommissionär Barnier att han i mig har en allierad som agerar för den här idén , som jag anser vara generös och europeisk .
Herr talman , herr kommissionär , kära kolleger !
Jämfört med hur ofta det uppträder stormar i andra områden i världen , är vi i Europa relativt förskonade .
Trots detta har stormarna under den sista decemberveckan visat vilka följder de kan få , och att vi också kommer att få stora problem .
Alla som åkte till Strasbourg med bil eller järnväg kunde övertyga sig om hur stormen rasat också i Alsace .
Jag vill därför uttala min medkänsla med alla medborgare i de regioner där stormen rasade så vilt , och samtidigt här i kammaren påpeka vikten av att stödja regionerna och människorna .
Vi alla vet att det i morgon lika gärna kan vara en annan region i Europa som drabbas på liknande sätt .
Det gäller nu att så snabbt som möjligt ta till vara dessa vindfällen .
Ty var och en vet att vi kan drabbas av ännu större katastrofer , om vindfällena får ligga kvar för länge i skogen .
Det måste också påpekas att exempelvis barkborren finner den bästa grogrunden för sin utbredning och för sina larver i vindfällena , och att det därigenom orsakas följdskador , som vi i dag ännu inte kan få någon uppfattning om .
Därför är det absolut nödvändigt att ta till vara vindfällena redan innan den varma årstiden börjar .
Den verkliga omfattningen av skadorna inom skogsbruket kommer vi att få reda på först om tiotals år .
Ty vi vet alla hur lång tid ett träd behöver på sig för att växa .
Här räknar man i årtionden , och inte i år .
Dessutom vill jag påpeka att det inom skogsbruket säkert inte bara gäller träproduktion , utan att de skyddade och de skyddande skogarna är en väsentlig faktor i vissa regioner .
Jag vill därför med stolthet säga att de österrikiska utbildade skogsarbetarna också är beredda att ...
( Talmannen avbröt talaren . )
Herr talman !
Vår djupaste medkänsla går till alla dem som drabbades av stormarna .
Ibland är vi inom gemenskapen egentligen inte medvetna om vad som händer i andra länder .
I Irland var mediatäckningen av det sjunkna tankfartyget väldigt liten .
Jag ombads berätta om konsekvenserna av stormarna i Irland .
Vi hade stark vind och ett långvarigt skyfall utan motstycke som lades till de svårigheter som redan fanns och resulterade i att hundratals hektar översvämmades och ibland lades under så mycket som 45 centimeter vatten .
Vi upplevde den mänskliga misären med översvämmade hem och gårdar , utan hälsovård och dricksvatten , och de miljömässiga katastroferna med E-kolibakteriesmittat vatten .
Jag talade med jordbrukare vars tackor fick missfall efter att ha druckit av det infekterade vattnet .
Naturliga livsmiljöer förstördes .
Därför ber jag er komma ihåg Irland i detta speciella fall .
Jag tackar kommissionären och stöder honom mycket starkt vad gäller hans europeiska insatsstyrka .
Herr talman , herr kommissionär , mina damer och herrar !
Jag ansluter mig till alla dem som har uttalat sin solidaritet med offren för stormen .
Jag vill också än en gång peka på betydelsen för skogsbruket i hela Europa .
Ty vi kommer ju att i alla områden i Europa få massiva effekter på skogsbruket , och jag tror att man här långsiktigt måste överväga hur man skall hantera sådana problem i framtiden .
Vi vill säkert inte ha någon organisation av marknaden för skogarna , men vi måste eventuellt skapa ett system , kanske även i samarbete med de privata försäkringsbolagen , och tillsammans med dem på något vis mildra sådana effekter för dem som drabbats .
Vi kommer tyvärr även i framtiden att tvingas räkna med dylika svåra katastrofer .
Det finns sådant som tyder på det , det har redan berörts här , det finns inga bevis , men tecken som tyder på att det ökande antalet stormar över hela världen har att göra med miljökastastrofen .
Forskarna är naturligtvis ännu inte eniga .
Men de flesta är relativt säkra på att om vi fortsätter med utsläppet av växthusgaserna så kommer dessa stormar naturligtvis att drabba oss ännu hårdare i det århundrade som just har börjat .
Jag tror att vi än en gång bör erinra om ett förslag som väcktes av en tidigare kollega till oss , Tom Spencer , här i kammaren ; enligt det bör vi inte ge stormarna några kvinnliga eller manliga förnamn , utan döpa dem efter dem som orsakar växthuseffekten - han nämnde då oljekoncernerna .
Här bör man dock säkerligen undanta Shell och BP , eftersom de har ändrat sin politik och inte bara satsar på försäljning av miljöskadliga fossila bränslen , utan också investerar i framtidsdugliga energiformer .
Detta sammanhang måste vi inse ; jag håller inte med dem som schablonmässigt säger att växthuseffekten bär skulden för denna storm , men att vi måste befara ytterligare katastrofer , om vi inte snabbt växlar spår , det är relativt säkert !
Herr talman !
Först skulle jag vilja tacka er för att ni förlängde debatten så att den blev sammanhängande .
Sedan skulle jag vilja säga att jag , i egenskap av kommissionär men också som fransk medborgare , blev oerhört rörd av de bevis på sympati och solidaritet som uttrycktes av många parlamentsledamöter från hela unionen .
Tack vare debatten gav de en aning om det jag tror på : ett Europa som inte kan sammanfattas som en stormarknad , utan ett Europa som också är mänskligt .
Jag skulle vilja tacka Scallon , Martin , McCartin , González Álvarez och Savary , som i synnerhet anammade och stödde den idé som jag försvarar , nämligen en lösning som i högre grad betonar det gemensamma , det praktiska genomförandet och tydlighet när det gäller civil säkerhet och civilt skydd , vilket skulle kunna ta sig uttryck i en europeisk civil säkerhetsstyrka .
Vi kommer att fortsätta att arbeta med den idén och rapportera för er under den närmaste tiden .
Många bland er - och jag har uppmärksamt lyssnat till Gebhardt , Patrie , Isler Béguin , Souchet , Gollnisch , Savary - sade att det inte finns tillräckligt med pengar , eller snarare att det inte finns ytterligare pengar .
Men , mina damer och herrar ledamöter - jag har varit parlamentsledamot under en mycket lång tid , så jag skall inte undervisa er - ni kan budgeten , ni känner till de allmänna bestämmelserna för strukturfonderna ; ni röstar igenom budgeten och ni vet alltså mycket väl inom vilka ramar jag arbetar .
Jag vill inte berätta sagor , jag vill göra ett seriöst arbete .
Detta hindrar mig inte från att tycka att man faktiskt skulle kunna återupprätta budgetposten om katastrofhjälp , med strikta ramar och med en ytterst detaljerad kravspecifikation , även om den posten endast avsåg några miljoner euro .
En summa som saknar samband med vidden av de katastrofer och deras konsekvenser som vi nu genomlider .
Ni känner till budgeten .
Det är inom den ramen jag arbetar , och vad gäller mitt eget ansvarsområde försöker jag att tillsammans med Diamantopoulou , för mål 3-budgeten , och Fischler , för Europeiska utvecklings- och garantifonden för jordbruket ( ( EUGFJ ) , se till att vi bemöter katastroferna såväl omedelbart som på medellång sikt , och att vi därmed gör EU-pengarna så effektiva som möjligt .
Jag motsätter mig således inte att budgetreglerna utvecklas , det kommer vi att tala om igen inför nästa budget - kanske för att återupprätta katastrofposten som avskaffades för två år sedan , åtminstone på ett symboliskt plan .
I väntan på detta finns det mycket pengar , mycket pengar , och , herr Gollnisch , jag kan inte låta er säga att de är tillgängliga för en hypotetisk och avlägsen period .
De här pengarna finns att tillgå nu , det här året .
Och om de nationella myndigheterna gör sitt arbete , vilket jag tror att de gör , kommer dessa medel att kunna uppbådas för specifika problem och projekt redan i mitten av år 2000 och för de kommande åren .
Och pengar finns det i överflöd , även om de , i fråga om mål 2 , inte täcker alla olycksdrabbade områden .
I synnerhet dessa pengar kan uppbringas , och det säger jag till Liese och Mathieu - fru Mathieu , jag har inte talat om en skogspolitik som ligger i sin linda - och till Keppelhoff och Schierhuber .
När det gäller skogsbruket och återställandet av skogrikedomarna - något mycket viktigt för mig - finns det vid sidan av mål 2 möjligheter att oavsett områdesindelningen utnyttja de avsevärda medel som finns i EUGFJ , garantisektionen .
Jag skulle till sist vilja säga , eller upprepa , att alla dessa katastrofer inte behöver vara naturkatastrofer .
Det säger jag med stor ödmjukhet .
Bland er finns ledamöter som är ytterst kompetenta och kunniga i dessa ämnen , även om jag tidigare har skrivit flera arbeten om ekologi och miljö .
Jag tror faktiskt att det finns katastrofer vilkas konsekvenser man skulle kunna begränsa med politisk vilja .
Jag tänker då på översvämningarna , men även stormarna .
Kronberger , Messner och González Álvarez tog upp de stora klimatfrågorna , och jag kan säga att det någonstans förmodligen finns en koppling mellan konsekvenserna av dessa naturkatastrofer och den förda politiken , där Europa måste bli en drivande och förebyggande kraft i viktiga miljöfrågor .
Herr talman !
Jag vill tacka er , och tacka parlamentet för att ha gett kommissionen tillfälle att uttala sig .
Nu kommer vi att arbeta , inom ramen för gällande budget och regler , för att se till att de medel som ni har ställt till vårt förfogande används på bästa möjliga sätt och så snabbt som möjligt , så att vi skall kunna hantera konsekvenserna av dessa katastrofer och ge ett ekonomiskt , politiskt och mänskligt svar till de familjer som har blivit allvarligt drabbade .
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum på torsdag .
 
Livsmedelssäkerhet Jag har erhållit sju resolutionsförslag som lagts fram i enlighet med artikel 37.2 i arbetsordningen .
Nästa punkt på föredragningslistan är meddelande om livsmedelssäkerhet och uttalande av kommissionen . .
Herr talman !
Det gläder mig mycket att kunna ta detta första tillfälle i akt att tillsammans med min kollega Liikanen för parlamentet dra upp huvudlinjerna i kommissionens vitbok om livsmedelssäkerhet , som antogs i onsdags , 12 januari .
Vid min utfrågning i september lovade jag att denna vitbok skulle levereras snabbt .
Jag är glad att vi har kunnat leverera den så snabbt .
Mellan tre och fyra månaders intensivt arbete sedan den nya kommissionen utsågs i september ligger till grund för vitboken .
Den bygger på de omfattande rådslag som har förekommit under de senaste åren sedan kommissionens grönbok om livsmedelslagstiftning utkom .
Den avspeglar också våra erfarenheter från nyligen aktuella larmrapporter om sådant som dioxin och slam liksom från BSE-krisen .
Vitboken avspeglar också detta parlaments intressen , vilka ni har beskrivit både för ordförande Prodi och för mig vid de många tillfällen då vi har debatterat livsmedelssäkerhet i denna kammare sedan kommissionen utsågs .
Jag behöver inte påminna er om att konsumenternas förtroende för Europas livsmedelssäkerhetssystem allvarligt har påverkats av kriser och larmrapporter under de senaste åren och månaderna .
Kommissionen har förbundit sig att återskapa detta förtroende genom att skapa världens mest moderna och effektiva system för livsmedelssäkerhet .
När jag lanserade vitboken förra veckan sade jag att kundvagnen är ett av de mest kraftfulla vapnen på denna jord .
Europas konsumenter fattar de mest omdömesgilla besluten .
Om deras förtroende rubbas avspeglar inköpsbesluten detta .
Detta har i sin tur dramatiska konsekvenser för jordbrukare , producenter och industrin i allmänhet .
I en bransch som omsätter omkring 600 biljoner om året kan även en liten nedgång i förtroendet få betydande konsekvenser .
Inom den agrara livsmedelssektorn och jordbrukssektorn finns över 10 miljoner anställda .
Ett högt förtroende är en förutsättning för att öka sysselsättningen och konkurrenskraften .
Denna förtroendekris har också fått den olyckliga men oundvikliga konsekvensen att konsumenternas förtroende för system och institutioner på nationell och europeisk nivå som skall övervaka och säkerställa högsta möjliga livsmedelssäkerhet har försvunnit .
När jag säger allt detta vill jag också slå fast att Europa trots detta har en av världens bästa livsmedelsindustrier och också ett av de säkraste systemen för livsmedelskontroll .
Utmaningen är att göra systemet till de allra bästa .
Det övergripande syftet med vitboken om livsmedelssäkerhet är därför att skapa erforderlig lagstiftning och strukturer som kan garantera konsumenterna högsta möjliga hälsoskydd vid livsmedelskonsumtion .
Vi sätter upp en krävande och ambitiös dagordning för förändring .
Kommissionen kommer att behöva parlamentets fulla stöd om vi skall kunna uppnå våra mål enligt tidsplanen .
Vi kommer också att behöva rådets och andra nyckelfunktioners fullaste stöd .
I vitboken om livsmedelssäkerhet beskrivs en omfattande uppsättning åtgärder som fordras för att komplettera och modernisera dagens livsmedelslagstiftning inom EU .
Alla dessa åtgärder syftar till att göra den mer konsekvent , begriplig och flexibel .
Vi vill verka för en bättre tillämpning av denna lagstiftning och ge konsumenterna större öppenhet .
I den detaljerade handlingsplanen om livsmedelssäkerhet i vitboken finns en preciserad tidtabell för åtgärderna under de närmaste tre åren .
Över 80 åtgärder planeras .
Vårt mål är att ha skapat en konsekvent och modern livsmedelslagstiftning vid utgången av år 2002 .
Vi planerar också att etablera en europeisk livsmedelsmyndighet år 2002 , som ett viktigt komplement till den nya livsmedelssäkerhetslagstiftningen .
Denna idé kommer att bli föremål för mycken analys och debatt .
Den har redan gett upphov till många kommentarer , inklusive reaktioner från parlamentsledamöter .
Det kapitel i vitboken som handlar om att skapa en europeisk livsmedelsmyndighet är klart utformat för att locka fram åsikter och kommentarer .
Vi vill ha in synpunkter på våra planer före slutet av april .
Jag kommer att återkomma till detta rådslag om några ögonblick .
Kommissionen anser att det krävs en övergripande strukturell förändring av vårt system för livsmedelssäkerhet för att säkerställa de nära besläktade målen att garantera högsta livsmedelssäkerhet och återställa konsumenternas förtroende .
Varför skulle en europeisk livsmedelsmyndighet vara en viktig del av denna förändring ?
Den första nyckelfrågan är oberoende .
Huvudaktörerna , däribland konsumenterna , söker ett system som är oberoende och som upplevs som fristående från alla lagstadgade intressen .
Vi måste också garantera förträfflighet och öppenhet .
Vi har gjort många framsteg under de år som har gått sedan det reformerade systemet med vetenskapliga råd antogs som en konsekvens av BSE-krisen .
Emellertid menar kommissionen att vi måste gå längre .
Vi måste skapa ett permanent och verkligt oberoende , utmärkt och öppet system för riskvärdering .
Myndighetens huvuduppgift kommer att vara riskvärdering inom livsmedelssäkerhetsområdet .
Vi tänker oss att de uppgifter de befintliga fem vetenskapliga kommittéerna som sysslar med livsmedelssäkerhet har skall överföras till myndigheten .
De kanske inte överflyttas med sin nuvarande form eller struktur - detta är en fråga som vi vill ha synpunkter på innan vi framlägger våra slutliga förslag om att inrätta myndigheten .
Om vi emellertid bara skulle föreslå en ommöblering skulle detta naturligtvis inte vara tillräckligt .
Som klargörs i vitboken måste den nya myndigheten ge ett mervärde .
Jag anser att det nuvarande systemet med vetenskapliga råd behöver förstärkas .
Inom denna myndighet tänker jag mig ett mycket starkare vetenskapligt och annat stöd för de oberoende vetenskapsmännen .
Jag förställer mig också att myndigheten kommer att vara mycket mer förebyggande än vårt nuvarande system - att förekomma snarare än reagera , att identifiera frågor innan de blir till kriser .
Detta förebyggande tillvägagångssätt bör bli myndighetens ledstjärna .
För att myndigheten skall kunna förebygga identifieras i vitboken ett antal nya områden som den skulle hantera .
Här ingår en omfattande informationsinsamling och övervakning , samordning av vetenskaplig information inom EU och uppbyggande av starka nätverk med livsmedelssäkerhetsenheter och -organ i medlemsstaterna .
Vi tänker oss också att myndighetens befogenheter skall omfatta driften av ett utbyggt snabbvarningssystem för problem med livsmedel och foder .
Kommissionen har beslutat att det varken är lämpligt eller möjligt att överlåta riskhantering till myndigheten .
Vi anser att beslut som gäller riskhantering fortfarande skall förbehållas kommissionen , parlamentet och rådet .
Jag ber inte om ursäkt för denna inställning för jag är övertygad om att den är riktig .
Naturligtvis finns det de som skulle hävda att vi bör ge en sådan myndighet lagstiftande makt .
Jag accepterar inte detta synsätt och tillbakavisar det med viss hetta .
Så sent som förra året ändrades fördraget så att parlamentet fick en mycket större roll i lagstiftningsprocessen .
Att i detta skede ge en myndighet denna roll vore enligt min mening ett steg tillbaka och skulle innebära en urvattning av det demokratiska ansvaret .
Jag är mycket intresserad av att höra parlamentets synpunkter i denna fråga .
Det finns också de som hävdar att kommissionen egentligen skulle kunna ignorera den nya myndighetens råd .
Jag tillbakavisar även detta resonemang .
Hur kan en kommissionär för hälsa och konsumentskydd avslå eller ignorera välgrundade vetenskapliga råd från oberoende källor om livsmedelssäkerhet ?
Skulle detta ligga i Europas medborgares intresse ?
Enligt min åsikt skulle de flesta definitivt inte göra det , om inte ett sådant tillbakavisande av de vetenskapliga argumenten hade sunda skäl , kunde försvaras rationellt och var helt rättfärdigat .
Det är svårt att tänka sig en sådan situation .
Jag kan försäkra er här i dag att kommissionen kommer att ta full hänsyn till myndighetens vetenskapliga råd när den utövar sin riskhanteringsfunktion .
Jag har redan sagt att myndigheten kommer att ansvara för att utveckla nätverk med nationella livsmedelssäkerhetsenheter och -organ i medlemsstaterna .
Detta är en stor uppgift .
Vi måste utveckla en större säkerhet i den vetenskap som bär upp livsmedelssäkerheten i Europeiska unionen .
Myndigheten måste bli en auktoritet för vetenskaplig rådgivning och information om livsmedelssäkerhet .
Denna situation skapas inte genom myndighetens blotta tillkomst utan kommer att framträda efter hand i takt med att självförtroendet stiger inom myndigheten själv .
Jag tror inte att vi kan vara föreskrivande gentemot vetenskapen och råd som grundas på vetenskap .
I och med att dynamiska nätverk utvecklas med nationella livsmedelssäkerhetsenheter och -organ kommer dock myndigheten att bli dominerande på den europeiska scenen .
Jag vill också gärna höra parlamentets synpunkter på detta .
Som en integrerad del i en mervärdesstruktur föreslås i vitboken att myndigheten skall ha en huvudroll inom riskkommunikation : att sprida komplicerad vetenskaplig information på ett konsumenttillvänt sätt , att vara den självklara och oundgängliga instans man vänder sig till för de allra senaste riskuppgifterna , att vara mycket synlig , att berätta goda nyheter om livsmedel , att vara förebyggande .
Vitboken innehåller också mycket viktiga förslag vad kontrollen beträffar .
Detta är en enormt viktig beståndsdel i systemet av avprickning och avrapportering för att tillse att medlemsstaterna och aktörerna uppfyller gemenskapens lagstiftning .
Jag vill se en riktig inre marknad i funktion på kontrollområdet .
I detta sammanhang föreslår vi också att den kontrollfunktion som utövas av kontoret för livsmedels- och veterinärfrågor i Dublin stärks betydligt .
Denna reviderade gemenskapskonstruktion skulle ha tre grundstenar : operativa kriterier som fastslås på gemenskapsnivå , riktlinjer för gemenskapskontroll och ett ökat administrativt samarbete för att utveckla och bedriva kontroll .
Som en del av våra förslag på detta område - som jag har för avsikt att lägga fram mot slutet av året - kommer jag att granska om kommissionen behöver ges ytterligare maktmedel som komplement till förfaranden vid överträdelser .
Dessa skulle kunna inkludera att innehålla finansiellt stöd från gemenskapen eller att återkräva medel som redan överlämnats till en medlemsstat .
Dessa förslag skall ses som en del i vår strävan att ha världens strängaste normer för livsmedelssäkerhet , öka konsumenternas förtroende och vidga marknaderna för jordbrukare och producenter i unionen .
Förutom förslagen om en ny europeisk livsmedelsmyndighet och ett förstärkt kontrollsystem på gemenskapsnivå innehåller vitboken förslag till en handlingsplan med ett brett spektrum åtgärder för att förbättra gemenskapens lagstiftning och göra den mer konsekvent , vilka täcker alla aspekter av livsmedelsprodukter från bondgården till köksbordet .
Här beskrivs över 80 enskilda åtgärder som planeras under den period vi har framför oss i syfte att täppa till de identifierade kryphålen i dagens lagstiftning .
Den nya rättsliga ramen kommer att omfatta djurfoder , djurens hälsa och välfärd , hygien , föroreningar och residuer , nya födoämnen , tillsatser , smakämnen , förpackning och bestrålning .
Den kommer att innehålla ett förslag till generell livsmedelslagstiftning som inbegriper principerna om livsmedelssäkerhet såsom fodertillverkares , jordbrukares och livsmedelshanterares ansvar , om att foder , livsmedel och ingredienser skall kunna spåras , om ordentlig riskanalys genom till exempel riskvärdering - det vill säga vetenskaplig rådgivning och informationsanalys - om riskhantering - det vill säga reglering och kontroll - riskkommunikation och tillämpning av försiktighetsprincipen om och när det är lämpligt .
Vad försiktighetsprincipen beträffar kan jag tillägga att kommissionen för närvarande håller på att slutföra ett meddelande som jag förväntar mig skall antas mycket snart .
Jag ser fram emot ett nyttigt utbyte av åsikter i eftermiddag med parlamentets ledamöter , som förstås skulle ha föredragit att göra detta förra veckan om något lämpligt parlamentsforum hade funnits tillgängligt .
Mot bakgrund av mina kontakter med ordförandena i berörda utskott inser jag emellertid att detta inte lät sig göras .
Men jag vet också att vi kommer att få många fler tillfällen att överväga förslagen om en myndighet i vitboken under de kommande månaderna .
Vi har nu ett antal månader på oss för att avhålla den nödvändiga debatten om kommissionens idéer om vitboken om inrättandet av en europeisk livsmedelsmyndighet .
Parlamentet kommer att spela en viktig roll i denna debatt .
Parlamentet spelade en avgörande roll i Europas svar på BSE-krisen .
Det har varit särskilt aktivt sedan dess för att sätta medborgarnas oro om livsmedelssäkerheten i förgrunden .
Jag väntar mig att parlamentets bidrag till debatten om myndigheten skall bli lika betydande och konstruktivt .
Även om vi har ett antal månader på oss till slutet av april för att debattera denna fråga och samla in våra synpunkter inser jag fullkomligt att detta också är en mycket stram tidtabell .
Jag skulle därför vilja be parlamentet att vidta lämpliga åtgärder för att tillse att dess åsikter formuleras så snabbt som möjligt .
Det är viktigt att kommissionen får dra nytta av parlamentets bidrag till formandet av det som är tänkt att bli en viktig del i arbetet för att föra upp skyddet av konsumenternas hälsa till ett nytt plan och därigenom återställa konsumenternas förtroende för Europeiska unionens politik för livsmedelssäkerhet .
Den europeiska livsmedelsmyndigheten kommer att bli en huvudaktör i EU : s politik för livsmedelssäkerhet under kommande år .
Det är viktigt att vi ger den rätt ingredienser .
Herr talman !
Jag tackar kommissionären för hans uttalande .
Jag skulle vilja uttrycka min uppskattning av den arbetsfördelning ni har gjort och av att livsmedelsfrågorna kommer att förbli en angelägenhet för de europeiska institutionerna , inklusive kommissionen och parlamentet .
Detta är alldeles rätt inställning .
Men det finns ett ord som jag inte har hört er nämna i kväll .
Jag hoppas att vi kan reda ut det här .
Vi behöver en livsmedelslagstiftning , som ni sade , och vi behöver komma överens om detta .
Det är väldigt viktigt att vi inbegriper ansvaret i denna process .
Det är detta ord jag menade .
Problemet hittills är att skattebetalarna har betalat när någonting har gått fel .
Detta kan inte fortgå .
När vi har en kris måste vi klart slå fast i förväg att om det finns ett problem är de som är upphov till det betalningsansvariga .
Herr talman !
Det var en mycket bra vitbok , det vill jag inte förneka .
Mina frågor gäller positivlistan för djurfoder .
Det är oklart i er vitbok .
Hur ser er tidsplan ut , hur snabbt kommer ni att lägga fram en positivlista ?
När kommer det att ställas samma krav på djurfoder och uppfödning som på tillverkning av livsmedel och kontroll av livsmedelstillverkningen ?
Den sista delen av min fråga : När kommer BSE-tester att bli obligatoriska i alla medlemsländer ?
Även där är ni , beträffande förpliktelsen , något oklar i er vitbok .
Tack för ert uttalande , herr kommissionär .
Jag anser att de linjer ni har dragit upp vad beträffar livsmedelssäkerhetsmyndigheten speglar verkligheten .
Medlemsstaterna skulle inte acceptera ett reglerande organ , så det är ingen större idé att ni föreslår ett .
För vissa delar av livsmedelsindustrin krävs uppenbarligen bättre lagstiftning och detta står klart i fråga om livsmedel och djurfoder .
I egenskap av ordförande i ett utskott som verkar komma att ägna sig nästan uteslutande åt livsmedel under de kommande tre åren måste jag dock fråga : om Europa har det säkraste systemet för kontroll av livsmedel , som ni sade , varför behöver vi då 24 nya direktiv och förordningar och 20 nya ändringsdirektiv ?
För det andra , kommer inte detta att förvärra problemet med för mycket reglering från Bryssel och för litet tillämpning i medlemsstaterna ?
Vi ser fram emot en givande dialog med er om detta .
Vad utvidgningen beträffar : vilka planer har kommissionen på att dra in ansökarländerna i debatter om dessa nya lagar , under förutsättning att kommissionen verkligen förväntar sig att de lagar som planeras i vitboken skall utgöra en del av gemenskapens regelverk senast år 2003 ?
Herr talman !
Först av allt skulle jag vilja tacka Ahern , Roth-Behrendt och Jackson för deras stöd för vitboken .
Det tycker jag är uppmuntrande och jag ser fram emot ytterligare diskussioner med dem och med andra parlamentsledamöter om de frågor de tog upp .
Ahern tog upp frågan om ansvar .
Detta tas naturligtvis inte upp särskilt i vitboken förutom hänvisningen till det faktum att vi kommer att skapa bestämmelser - och det finns redan några - om möjligheterna att spåra livsmedel .
När väl detta är gjort kan frågor som ansvar tas upp .
Jag har trots min bakgrund inte helt och i detalj övervägt frågor som sammanhänger med och omger ansvarsfrågorna , men jag tror att det mycket väl kan vara subsidiaritetsfrågor involverade .
Men jag har noterat ert förslag och kommer att överväga det ytterligare .
Roth-Behrendt frågade mig om upprättandet av en positiv lista .
Det är en av de frågor vi tar upp i bilagan till lagförslaget och avsikten är att upprätta en positiv lista för fodermaterial .
För närvarande är listan , som jag säger , en negativ lista som fylls på vid behov .
Upprättandet av den positiva listan är en av de frågor som behandlas i bilagan som har ett datum åsatt , år 2002 faktiskt .
Det snabba varningssystemet för foder är någonting vi har identifierat som en lucka i lagstiftningen .
Snabb varning finns för livsmedel men inte för foder .
Detta är olyckligt och det är fel , och vi tror att det är viktigt att påpeka det och införa lagstiftning som täpper till denna lucka , och detta skall göras .
Medlemsstaternas arbete med BSE och införandet av stickprovstest för att identifiera infektionsnivåer i medlemsstaterna pågår .
Jag vet att Roth-Behrendt har frågat mig om detta förut och jag sade att jag tyckte att det gick snabbt framåt , men jag har förstått att ärendet befinner sig på intern remiss i kommissionen och att arbete pågår .
Jag hoppas att jag nästa gång ni ställer frågan kommer att vara i stånd att ge er mer detaljerad information .
Jackson inriktade sig på det faktum att det finns 24 nya och 20 ändringsakter i lagstiftningen och frågar om detta innebär överreglering .
Jag skulle vilja säga att de rättsakter vi har skiljt ut syftar till att täppa till luckor i gällande lagstiftning .
Det handlar inte så mycket om att skapa nya system för ytterligare reglering , även om detta är en del av det , utan om att identifiera var det finns luckor och kryphål i kedjan från bondgård till middagsbord och täppa till dem .
Det finns en hänvisning till ansökarländerna och detta är någonting vi tänker på .
Normer för livsmedelssäkerhet och också andra säkerhetsfrågor är naturligtvis av avgörande betydelse för utvidgningen och detta är en fråga jag har tagit upp med Verheugen .
Herr kommissionär !
Vissa medlemsländers okunnighet har fört oss in i en stor livsmedelskris i Europa , och jag är , tyvärr , än en gång irriterad över att rådet i sin helhet återigen saknas i dag , när ni lägger fram detta intressanta meddelande .
Jag skulle gärna vilja höra av er hur ni skall se till att en sådan ny myndighet , vad den än må heta i detalj , även får inflytande på rådet , vem i denna myndighet som skall bestämma , och vem som skall dela ut uppdragen .
Naturligtvis får vi inte föreskriva något om innehållet , men jag insisterar redan på att parlamentet efter Maastricht och Amsterdam skall behålla sin rätt och rent av bygga ut den .
Jag är mycket oroad över att vi återigen kan få en myndighet , som flyger anonym som en satellit över Europa ; en sådan myndighet skulle jag älska lika mycket som djävulen älskar vigvattnet .
Jag hoppas att det inte kommer att ske !
Även jag välkomnar vitboken .
Men planerar ni att livsmedelssäkerhetsmyndigheten skall ha tillräcklig makt för att förhindra något liknande det köttkrig vi har haft och Frankrikes vägran att häva importförbudet ?
Ni nämnde att kommissionen har möjlighet att hålla inne anslag och bidrag för länder som agerar på det sätt som Frankrike agerar .
Skulle ni då också föreslå att kommissionen kan göra interimsbetalningar till exempel , liknande de brittiska jordbrukare ber om för närvarande ?
Herr talman , herr kommissionär !
Vid ett informationsmöte i förra veckan sade ni att EU : s livsmedelsmyndighet enligt er uppfattning inte borde förläggas på en avlägsen ort , men ni sade inte vad ni menade med denna avlägsna ort .
Den verksamhet som EU-enheten i Dublin bedriver har exempelvis visat att det geografiska avståndet i dag inte är något hinder för effektiv påverkan och kontakt .
Man har sagt att den kommande livsmedelsmyndighetens viktigaste uppgifter är att samla in , publicera och samordna data , utfärda rekommendationer i syfte att utveckla livsmedelssäkerheten och - som ni konstaterade - samla in vetenskapliga yttranden och göra informationen lättillgänglig och lättförståelig för konsumenterna .
Allt detta kan med hjälp av dagens teknik skötas var som helst inom Europeiska unionens område .
Jag frågar därför , vad grundar ni er uppfattning om lokaliseringen på ? .
( EN ) Vad beträffar myndighetens utformning : för det första kommer den att anställa egna vetenskapsmän som kommer att hålla kontakt med och rådfråga vetenskapsmän som är experter på de just de områden som för tillfället är aktuella .
Dessutom kommer livsmedelssäkerhetsmyndigheten att ha en styrelse .
Ni kommer att märka av vitboken att vi inte har gått in på detaljer om hur denna styrelse skall vara sammansatt .
Detta är en fråga som jag förväntar mig att parlamentet och kommissionen kommer att diskutera under de kommande veckorna och månaderna .
Jag föreställer mig att styrelsen kommer att bestå av finansiärerna eller av företrädare för dessa .
I det förslag jag skall lämna till kommissionen i september måste dess funktion beskrivas i detalj .
Vi har inte gjort det än , men det kommer att göras i september .
Jag väntar mig inte att styrelsen skall tala om för vetenskapsmännen hur de skall sköta sitt arbete .
Det skulle eliminera de vetenskapliga rådens oberoende .
Men den kommer att ha en generell befogenhet , särskilt till exempel för att kräva att myndigheten granskar vissa områden som behöver utforskas .
Florenz frågar om parlamentet kommer att ha någonting att säga till om här .
Det är en fråga att överväga och diskutera .
Det kan finnas ett antal åsikter om det .
Vissa kanske intar ståndpunkten att det vore olämpligt att parlamentet eller parlamentsledamöterna - eller rent av av parlamentet utsedda ledamöter - sitter med i styrelsen .
Andra kanske anser att det skulle vara en nyttig övning om parlamentet , via ombud eller ledamöterna själva , skulle få en möjlighet att diskutera vilka frågor som skall undersökas .
Det tål att tänka på , men det är inte uteslutet .
Florenz tog också upp frågan om anonymitet .
Jag är glad att han tog upp den eftersom det är särskilt viktigt att denna myndighet har en hög profil .
Den måste synas .
Den måste vara känd .
Konsumenterna i Europeiska unionen måste veta att livsmedelsmyndigheten finns .
Myndighetens VD bör vara någon som är känd , någon som kanske regelbundet medverkar i TV-program om livsmedelsfrågor , särskilt vad gäller de goda livsmedelsnyheterna om näringsvärden , kosthållning och liknande , så att konsumenterna känner till att en sådan myndighet finns om en ny livsmedelskris uppstår .
De skall vara medvetna om att de har hört talas om myndigheten tidigare under andra omständigheter och förhoppningsvis ha ett grundförtroende som redan har byggts upp genom myndighetens uttalanden .
Det är därför av avgörande betydelse att myndigheten inte är anonym .
Den måste synas .
Jag kommer att göra allt som står i min makt för att verka för att myndigheten får denna höga profil .
Lynne frågar om myndigheten kommer att ha tillräcklig makt .
Jag misstänker att frågan gäller var myndighetens befogenheter börjar och slutar och var livsmedelssäkerhetsmyndigheter i medlemsstaters ansvar och behörighet börjar och slutar .
Det skulle krävas en växelverkan på vetenskaplig nivå .
Det vore helt klart inte önskvärt med en situation där det uppstår motsättningar mellan vetenskapsmän som arbetar för eller är konsulter till livsmedelssäkerhetsmyndigheten på gemenskapsnivå och någon vetenskaplig åsikt på medlemsstatsnivå .
Detta är en icke önskvärd situation , en situation vi inte vill se i framtiden .
Det finns ett antal saker som undergräver konsumenternas förtroende , och informationsbrist är en av dem .
Men information som innehåller grundläggande meningsskiljaktigheter mellan vetenskapsmän i viktiga frågor som gäller livsmedelssäkerhet är också något som inger stor oro .
Vi måste försöka undvika detta och skapa strukturer som säkerställer att det finns ett ordentligt informationsutbyte mellan vetenskapsmännen , att rådslag och diskussioner genomförs till fullo och att myndigheten på gemenskapsnivå har möjlighet och mandat att fråga oberoende vetenskapsmän i alla medlemsstaterna och kanske rent av längre bort , när experter finns annorstädes , om råd och åsikter .
Med tiden kommer , som jag sade nyss , inte bara myndigheten att få en tydligare profil utan dess expertis , dess moraliska auktoritet , kommer att öka i takt med att tiden går så att dess åsikter accepteras och inte ifrågasätts .
Denna situation kan vi uppnå med tiden .
Man kan inte lagstifta fram konsumenternas förtroende .
Det är någonting man vinner med åren .
Kommissionen kommer emellertid att ha möjlighet att tillse att myndighetens åsikter i vetenskapliga frågor genomdrivs genom att lagstiftning antas , vilket är kommissionens , parlamentets och rådets funktion .
Jag inser att detta är en något tidsödande övning , men trots detta anser jag att införandet av lagstiftning som härrör ur myndighetens ståndpunkter är rätt väg att gå .
Om lagstiftningen inte följs kan detta hanteras i domstolarna på normalt sätt .
En av de frågor som vi kan komma att tvingas ta upp med tiden är frågan om svarstider under sådana omständigheter .
Jag tänkte se om någonting kan göras , så att vi får snabbare respons från domstolsprocessen .
Vad gäller anslag och bidrag : ja , vi har tagit hänsyn till denna fråga .
Den kommer att kräva juridisk rådgivning och detta kommer vi att begära , särskilt med tanke på att det kan ge ett snabbt svar på underlåtenhet att uppfylla gemenskapslag i avvaktan på ett domstolsutslag .
Vad gäller Lynnes fråga om interimsbetalningar : detta är en fråga som mycket väl kan tas upp i parlamentet , eftersom den gäller budgetfrågor .
Myller frågade sedan om myndighetens placering .
Inget beslut har fattats om detta annat än att säga att det är mer troligt att myndigheten placeras centralt än perifert .
Jag inser att FEO är placerat i Dublin och , trots att jag själv kommer från den delen av världen , måste jag acceptera att det inte är Europas centrum !
Men FEO befinner sig i en helt annan situation än livsmedelssäkerhetsmyndigheten .
FEO består av oberoende vetenskapsmän och veterinärer och så vidare som reser från någon plats där det finns en flygplats - och det har vi helt klart i Dublin .
Livsmedelssäkerhetsmyndigheten har en helt annan situation .
Den måste finnas nära kommissionen till följd av behovet av samverkan mellan de vetenskapsmän som arbetar för livsmedelssäkerhetsmyndigheten och de av oss som är involverade i lagstiftningsinitiativ .
En viktig del av kommunikationen mellan de två institutionerna kommer självfallet att bli att tillse att de av oss som sysslar med att göra upp lagförslag tydligt och klart förstår vad vetenskapsmännen menar , vilka problem de har identifierat , vilken lagstiftning som krävs för att ta itu med de frågor de tar upp .
På samma sätt kommer vetenskapsmännen att vilja ha något inflytande på utformningen av politik och lagstiftning för att tillse att lagstiftningen botar det onda de har identifierat .
Jag tycker det verkar önskvärt att en sådan myndighet är centralt placerad .
Vetenskapsmännen kommer att vara fast anställda , men det kommer också att bli nödvändigt att arbeta med vetenskapsmän på konsultbasis och under dessa omständigheter är det förmodligen bättre att de , eftersom de måste resa , förflyttar sig till en central plats , där återigen parlamentets strukturer och kommissionen och rådet är baserade .
Detta är min bedömning för tillfället .
Det kan bli ämnet för diskussion här och annorstädes och jag kommer att lyssna på alla förslag som framläggs , men min preliminära slutsats är att denna myndighet hellre bör vara centralt placerad än i periferin .
Jag befinner mig i en mycket svår position för jag kan inte ändra föredragningslistan .
Jag skulle vilja föreslå att ni tar upp detta med era politiska grupper och på talmanskonferensen .
Om ni känner att dessa sessioner efter ett uttalande från kommissionen är viktiga skulle jag föreslå att vi kräver mer tid än den halvtimme som är avsatt för dem .
Vid detta tillfälle har vi haft sex minuter frågor från ledamöterna och 29 minuter svar från kommissionären , samt hans uttalande .
Som ni ser är en halvtimme egentligen inte i närheten av vad som vore tillräckligt för en sådan sittning .
Jag hoppas att ni diskuterar detta i era politiska grupper så att vi kan få en mer välstrukturerad sittning med kommissionen vid framtida tillfällen .
Jag förklarar debatten avslutad .
 
Frågestund ( kommissionen ) Nästa punkt på föredragningslistan är frågor till kommissionen ( B5-0003 / 2000 ) .
Jag vill meddela att frågestunden kommer att pågå i cirka en timme och femton minuter .
Vi kommer dock att begränsa tiden något , eftersom tolkarna arbetar oavbrutet under dagens sammanträde .
Jag överlämnar ordet till Purvis för en ordningsfråga .
Jag protesterar mot att vi drar ned på tiden för frågestunden .
Det är ett av de få tillfällen då vanliga ledamöter har en chans att få tala och jag ber er att utöka den till en och en halv timme som på föredragningslistan .
Så säger föredragningslistan och jag anser att vi skall hålla oss till den .
Faktum är , käre kollega , att vi enligt föredragningslistan borde börja kl .
17.30 , och ni har klockan framför er .
Jag hoppas åtminstone att sammanträdet inte fortsätter långt in på natten .
Första delen Fråga nr 28 från ( H-0781 / 99 ) : Angående : Anläggning av kärnkraftverk i det jordbävningsdrabbade Turkiet De två senaste jordbävningarna i Turkiet som båda mätte över 7 grader på Richterskalan föder stor undran över att turkarna envist framhärdar med att uppföra dyra kärnkraftsreaktorer i Akköy - samtidigt som energiförråden från Ataturk-dammarna exporteras till tredje länder och EU gör nedskärningar i sin budget för att kunna bevilja pengar för restaureringsarbetena med anledning av de skador som jordbävningarna förorsakat .
De turkiska planerna för utvecklande av kärnkraft , som inte verkar ta hänsyn vare sig till de faror som dessa innebär för invånare eller ekosystem i Turkiet och angränsande områden , föder misstankar om att det kanske bakom dessa planer döljer sig medvetna beslut , som fattats av de turkiska politiska och militära makthavarna , om att tillägna sig kärnteknik som i framtiden skall möjliggöra framställning av kärnvapen .
Fog för dessa misstankar finner man bland annat i det faktum att landet har för avsikt att skaffa sig reaktorer av kanadensisk typ , det vill säga likadana som de reaktorer som finns i Indien och Pakistan .
Vilka åtgärder tänker kommissionen vidta för att kärnkraftsolyckor skall kunna undvikas och spridande av kärnvapen skall kunna hindras i ett land som önskar ansluta sig till EU och som spenderar enorma summor på program för utvecklande av kärnteknik samtidigt som det slukar europeiska medel beviljade av EU , medel som det erhåller i form av ekonomiskt bistånd ?
Jag överlämnar ordet till Verheugen som företrädare för kommissionen . .
( EN ) Kommissionen följer med intresse det planerade bygget av ett kärnkraftsverk i Akkuyu i Turkiet och inser vikten av att säkerställa att det nya verkets konstruktion följer högsta internationellt godkända standard för kärnenergisäkerhet .
Enligt vad vi har erfarit har inte beslutet om val av entreprenör tagits ännu .
Kommissionen noterar det faktum att Turkiet har undertecknat och ratificerat konventionen om kärnenergisäkerhet och att ansvaret för att bevilja tillstånd och reglera förläggning , konstruktion , igångkörning , drift och nedstängning av kärnkraftverk i Turkiet helt åvilar den turkiska atomenergimyndigheten .
Kommissionen har inget mandat att sätta upp gränser för beslut som fattas av något land om energiproduktion , kärnkraften inbegripen .
Som kommissionär Wallström berättade under utfrågningen i Europaparlamentet i september 1999 kommer kommissionen att ta upp frågan om kärnenergisäkerhet och strålskydd vid alla relevanta möten med den turkiska regeringen i framtiden och det gläder mig att kunna informera er om att jag kommer att ha ett möte med den turkiske utrikesministern om några dagar och förstås kommer att ta upp frågan .
Kommissionen är särkilt medveten om allmänhetens oro för den uppmätta seismiska aktiviteten i området kring Ecemis-förkastningslinjen i närheten av den plats där verket föreslås bli placerat .
Enligt information från Internationella atomenergiorganet tar man i verkets utformning hänsyn till möjligheten av jordbävningar som är kraftigare än några som någonsin har registrerats i området och mer än tio gånger kraftigare än den som uppmättes i Adana i juni 1998 .
Stora utformningsmässiga marginaler skapas för att säkerställa att verket kan drivas säkert i enlighet med miljöförhållandena på platsen .
Kommissionen är också medveten om oron för den möjliga avsikten att använda verket för att producera material till vapen .
Den noterar det faktum att Turkiet har undertecknat och ratificerat fördraget om icke spridning av kärnvapen och därefter har slutit ett omfattande avtal om garantier med Internationella atomenergiorganet .
Jag tackar för svaret .
Jag vill göra följande påpekande : Turkiet är nu kandidatland .
Genom detta projekt vill landet öka sin energikapacitet med 2 procent .
Samtidigt vill det förvärva reaktorer av typ Cadou från Canada , reaktorer som redan har använts för att framställa Pakistans och Indiens kärnvapen , som det har framkommit .
Mot denna bakgrund finns det en mycket allvarlig risk att någon vettvilling kommer fram till att den geostrategiska balansen i Kaukasus kräver att det i närheten finns ett land med kärnvapenteknik Detta är den politiska aspekten .
Jag övergår nu till den tekniska aspekten .
Säkerhetskoefficienten vid anläggningar av detta slag - och jag talar nu som ingenjör - har inget samband med att risken för reaktorhaveri ökar 10 eller 20 gånger .
När det råder tveksamhet , använder man i dessa fall simulatorer .
Vi kan emellertid inte använda simulatorer , när det gäller kärnkraft .
Därför måste alla områden med hög seismisk risk a priori vara uteslutna , när det gäller kärnkraftsanläggningar av denna typ .
Eftersom Europeiska unionen och kommissionen nu har andra möjligheter i fråga om Turkiet , bör man också diskutera vissa frågor som gäller säkerheten i området som helhet , men också frågan om Turkiets fredliga utveckling i Europeiska unionens sammanhang . .
( EN ) För några veckor sedan hade vi en debatt i parlamentet om kärnenergiäkerhet med speciell inriktning på kandidatländerna .
Jag har förklarat kommissionens inställning .
Man måste acceptera det faktum att det inte finns något regelverk i gemenskapen för kärnenergisäkerhet .
Så det vi gjorde var att använda politiska medel för att övertyga vissa kandidatländer om att vi måste ha nedstängningsplaner för somliga reaktorer som inte anses möjliga att uppgradera .
I fråga om Turkiet är det annorlunda .
Kärnkraftverket finns inte än .
Jag har redan sagt att Turkiet har undertecknat icke-spridningsavtalet och konventionen om kärnenergisäkerhet .
Om vi under fullbordandet av detta kärnkraftverk finner att det finns säkerhetsproblem kommer vi att diskutera detta med Turkiet .
Om slutsatsen är att Turkiet planerar att bygga ett kärnkraftverk som inte uppfyller normala europeiska säkerthetsnormer kommer vi att göra samma sak som med Litauen , Slovakien och Bulgarien .
Herr talman !
Kommissionären sade att Turkiet har undertecknat icke-spridningsavtalet och kärnenergisäkerhetsfördragen : varför skulle det finnas något som helst tvivel på att Turkiets kärnkraftverk inte skulle bli precis lika säkert som något annat i gemenskapen , och skulle kommissionären vara beredd att inta en något mer kraftfull ståndpunkt mot Souladakis i denna fråga ? .
( EN ) Jag anser att en parlamentsledamot har rätt att ta upp det han oroar sig och är rädd för .
Jag är inte orolig för detta .
Jag tror att Turkiet till fullo godtar normerna och kriterierna i konventionen om kärnenergisäkerhet och i icke-spridningsavtalet , men det finns otvivelaktigt en oro bland allmänheten i Europa och jag tycker att det är helt rätt att diskutera den här i parlamentet .
Fråga nr 29 från ( H-0786 / 99 ) : Angående : Vapen med utarmat uran Har kommissionen gjort några utredningar av hur staterna inom EU kan komma att påverkas av gränsöverskridande föroreningar som uppstått till följd av att det i Kosovokonflikten använts vapen med utarmat uran ?
Om inte : varför inte ?
Härmed överlämnar jag ordet till Wallström , som företrädare för kommissionen . .
( EN ) Tack för er fråga , herr Bowe .
Europeiska kommissionen har övervakat konfliktens miljökonsekvenser från det att Natoaktionen inleddes .
Redan i juni förra året finansierade kommissionen en första utredning .
Den genomfördes av det regionala utvecklingscentrumet för Central- och Östeuropa och slutsatsen var att ingen storskalig ekologisk katastrof hade ägt rum .
Denna första bedömning har inte ändrats av senare bevis eller analyser .
Kommissionen har också varit intimt inblandad i framtagandet av den rapport som nyligen utgavs av Förenta Nationernas miljöprogram - insatsstyrkan på Balkan .
Detta är den hittills mest detaljerade och omfattande rapporten om Kosovokrigets miljökonsekvenser och jag rekommenderar dem av er som ännu inte har tagit del av den att göra det .
Användningen av utarmade uranvapen var en av de många frågor som behandlades och denna rapport finns nu lätt tillgänglig , också på Internet .
Insatsstyrkan på Balkan hindrades av det faktum att det praktiskt taget inte fanns någon information om den faktiska användningen av dessa vapen under kriget .
På sin faktainsamlingsresa fann de inga tecken på kontamination i Kosovo .
Detta utesluter dock inte att områden i Kosovo kan vara kontaminerade med utarmat uranium .
Av en skrivbordsutvärdering tillsammans med en faktainsamlingsresa dras i rapporten slutsatsen att eventuella risker begränsas till ett område kring målet .
Framtida åtgärder kommer att genomföras inom ramen för stabilitetspakten för sydöstra Europa .
En särskild regional plan för rekonstruktion av miljön håller också på att tas fram .
Den kommer att bilda ramen för nödinsatser för att bekämpa krigsskador , om sådana skulle behövas .
Herr talman !
Först av allt ber jag att få tacka kommissionären för detta mycket matnyttiga svar .
Det är tydligt att kommissionen har övervägt detta problem , och jag är glad att man i de rapporter som hittills har framtagits granskar frågan ingående .
Men jag skulle vilja påpeka att oron för utarmade uranvapen gäller sättet de används på .
Detta uranium blir luftburet och man andas in det .
Det skulle nu faktiskt kunna vara så att delar av befolkningen i Kosovo bär på detta , med mycket mer långsiktiga effekter än man hittills kunnat fastställa .
Detta verkar vara det händelsemönster som har framkommit efter användningen av utarmade uranvapen i Gulfkriget .
Jag skulle därför vilja fråga kommissionen om den skulle vilja överväga att fortsätta övervakningen och under hur lång tid de skulle kunna tänka sig att i framtiden övervaka för att se vilka de långsiktiga konsekvenserna blir , inte bara av utarmade uranvapen utan också en del av de andra miljökonsekvenser vi vet har uppstått åtminstone lokalt i Kosovo ?
Hur länge kommer ni att fortsätta att utvärdera konsekvenserna av dessa vapen ? .
( EN ) Tack för den frågan , herr Bowe .
Vi måste återigen hävda att det fortfarande inte är bekräftat att utarmat uran användes i kriget och att inget utarmat uran har upptäckts under upprensningen i Kosovo .
Men de symptom och de problem ni nämnde kan finnas där , och de kan vara konsekvenser av användningen av utarmat uran .
Detta nämns också i rapporten .
Inga gränsöverskridande konsekvenser har upptäckts och de flesta vapnen måste ha använts inom Förbundsrepubliken Jugoslaviens territorium .
Problemet är att landets nuvarande politiska isolering innebär att tillträdet till detta område är begränsat .
Förenta nationerna har ett stort ansvar , för denna rapport vänder sig till dem , så de måste ta sitt ansvar .
Men genom denna regionala och miljömässiga rekonstruktionsplan kan vi fortsätta övervakningen och det bistånd vi kan ge och detta är , för närvarande , den slags ram vi kan använda för Europeiska unionens arbete .
Uppföljning är viktig och den ger medlemsstaterna , liksom Förenta nationerna och kommissionen , någonting att tänka på när den handlar om militära hemligheter och deras konsekvenser för miljön .
Den har också en långsiktig påverkan på tänkandet när det gäller användningen av detta slags vapen .
Herr talman , fru kommissionär !
Om några månader kommer återigen hundratusentals semesterfirare att fara till den adriatiska kusten och tillbringa sin sommarledighet där .
Som vi känner till från nyhetsrapporterna , har bomber och vapen fällts i närheten av kusten .
Kan ni bekräfta att semesterfirarna denna sommar kan bada riskfritt i Adriatiska havet , och har man planerat åtgärder för att undersöka hur hotbilden ser ut ? .
( EN ) Jag önskar att jag kunde garantera mycket , men tyvärr kan jag inte det .
Vi gör våra bedömningar utifrån rapporter som denna och de sändebud vi skickar ut för att kontrollera sådana här saker .
Det är detta vi grundar oss på när vi råder människor vad de skall göra .
Det vi har sett är att krig påverkar miljön på lång sikt och detta är farligt .
På miljöområdet har vi just antagit ett direktiv om föroreningar till havs .
Detta innefattar kulor och vapen och så vidare och är ett förvarningssystem .
Tyvärr kan vi inte utfärda garantier utan bara fortsätta att övervaka och försöka genomföra upprensningar .
Jag ville fråga kommissionären om det är sant att soldater från Natos väpnade styrkor som nu är stationerade i denna region genomgår särskilda kärnstrålningskontroller och att samma åtgärder inte tillämpas på civilbefolkningen i området ? .
( EN ) Jag kan inte svara på den frågan .
Jag har inte all den information som fordras för att svara ordentligt när det handlar om läkarkontroller och så vidare .
Vad vi vet från miljösidan är det jag redan har nämnt , att det nu finns en plan för rekonstruktion av miljön , men när det gäller läkarkontroller har jag ingen information .
Jag kan naturligtvis gå tillbaka och se om vi kan hitta den information som behövs .
Fråga nr 30 från ( H-0793 / 99 ) : Angående : Utnämning av ett särskilt EU-sändebud för Tibet För 1998 registrerade den tibetanska exilregeringen att över 4 000 tibetaner flytt över Himalayabergen till friheten med fara för liv och lem .
Många av flyktingarna drabbades därvid av allvarliga förfrysningsskador och många dog .
Den tvärpolitiska gruppen " Tibet " är mycket bekymrad över den allt värre situationen i Tibet och det står klart att Europeiska unionens nuvarande politik inte räcker till för att uppnå resultat vad gäller de svåra kränkningar av de mänskliga rättigheterna som tibetanerna i Tibet utsätts för varje dag .
Den tvärpolitiska gruppen " Tibet " , som verkligen oroar sig över de fortsatta kränkningarna av de mänskliga rättigheterna i Tibet och önskar stödja Dalai Lamas förslag om en dialog med den kinesiska regeringen för att lösa situationen i Tibet , uppmanar därför kommissionen att utnämna ett särskilt sändebud för Tibet , som skall sköta Europeiska unionens angelägenheter i denna fråga och bemöda sig om att föra samman tibetanska och kinesiska företrädare och / eller myndigheter i en dialog .
När kommer kommissionen att utnämna ett särskilt sändebud för Tibet ?
Jag överlämnar ordet till Patten , som företrädare för kommissionen . .
( EN ) Den oro Europaparlamentet uttrycker för Tibet delas av många .
Jag har länge trott på behovet att bestämt och rättframt för de kinesiska myndigheterna framhålla vår inställning i frågor om mänskliga rättigheter också i Tibet .
Europeiska unionen gjorde detta vid toppmötet mellan Europeiska unionen och Kina förra månaden och pressade kineserna i ett antal frågor om mänskliga rättigheter , däribland Tibet .
Vi uppmanade åter Kina att inleda en dialog med Dalai Lama .
Jag uppmanar igen Kina att göra det .
Vi kommer att fortsätta att ta upp Tibet med de kinesiska myndigheterna .
Vi gör också en del andra saker : inom dialogen mellan Europeiska unionen och Kina om mänskliga rättigheter har vi inriktat oss på ett antal praktiska steg , däribland att skicka ut experter på uppdrag till Tibet , planera program för utvecklingsbistånd och verksamhet inom hälsa och utbildning för tibetanerna .
Utnämningen av ett särskilt EU-sändebud för Tibet skulle främst vara en fråga för rådet att besluta om och parlamentet kanske vill ta upp frågan direkt med dem .
Men för egen del är jag inte säker på att det skulle bidra så mycket till våra ansträngningar i praktiken .
Det skulle troligen inte ha någon större inverkan på de kinesiska myndigheterna och vi har redan effektiva kommunikationskanaler med exiltibetanerna .
Jag tycker också att det är angeläget att akta sig för en exponentiell ökning av särskilda sändebud , hur gott syftet än är .
Herr talman , herr Patten !
Ni har naturligtvis utmärkta erfarenheter på grund av ni levt i Kina , och ni vet mycket väl hur tibetanerna anstränger sig för att åstadkomma en dialog , vilket hittills alltid har förhindrats .
Men om ert svar blir att vi skall vända oss till " Mister Gusp " , alltså till Solana , då befarar jag att det är en ensidig inriktning av utrikespolitiken .
Er ansats , som jag mycket väl rekommenderar som en sammanhållande ansats , har ju inspirerats av de mänskliga rättigheterna ; jag håller helt med om att vi måste ta oss an frågan om human rights .
Anhållandena , tortyren , stympningen av unga kvinnor och liknande , det är ju absolut diskussionsämnen som man kan ägna sig åt en hel kväll .
Om vi inskränker det och säger att rådet här också är ansvarigt , så befarar jag att dessa frågor om de mänskliga rättigheterna inte kommer i dagen tydligt nog .
Möjligheten att å ena sidan betona ekonomi och handel , men att mycket väl integrera de mänskliga rättigheterna , vore en åtgärd där vi egentligen satsar på kommissionens partnerskap , och inte säger att det är en fråga för rådet . .
( EN ) Låt mig klargöra för er vilken inställningen är .
Jag sade ingenting annat än sanningen när jag sade att utnämningen av särskilda sändebud är en fråga för rådet .
Det råkar vara så att vi hanterar de budgetmässiga konsekvenserna och rådet utser vederbörande .
Somliga kanske tycker att denna budgetfråga borde ses över på sikt .
Om vi lämnar det , för sådant är läget , innebär inte detta att vi inte har en åsikt och en befogenhet i fråga om mänskliga rättigheter , jag hoppas väldigt mycket att kommissionen under de närmaste månaderna kommer att kunna ta fram ett meddelande om mänskliga rättigheter där vi bland annat påpekar att det inte finns någon som helst motsättning mellan en omsorg om mänskliga rättigheter i Kina eller på andra håll i världen och Europeiska unionens handelsmässiga , kommersiella och andra intressen .
Jag har länge ansett att vi alla bör erkänna att de länder som det är bäst att göra affärer med är de länder som behandlar sina egna medborgare mest anständigt - överallt i världen .
Jag upprepar att vi har framfört vår uppfattning om Tibet till Kina .
Under de få månader som jag har varit kommissionär har det hänt två gånger , först i New York vid vårt möte med minister Tang och nyligen vid mötet i Peking och vi kommer att fortsätta att ge uttryck för denna oro .
Om jag får rekommendera en bok till er , eftersom jag inser att ni är intresserad av dessa frågor , rekommenderar jag en bok om Tibet som gavs ut precis innan jul och som är skriven av den framstående journalisten Isabel Hilton .
Herr talman !
Jag vill börja min tilläggsfråga med den tibetanska hälsningen , som betyder lycka och fred .
I Tibet handlar det inte bara om de mänskliga rättigheterna och miljön , utan det handlar om ett unikt kulturarv , som också kan förmedla viktiga värden till oss européer , exempelvis ro , stillhet , medkänsla , compassion , som Dalai Lama säger .
Frågan är nu vad kommissionen kan göra för att på ett mer konkret sätt stödja Hans Helighet Dalai Lama och hans förslag till en fredlig lösning av Tibet-frågan ?
Jag vill påpeka att om man inte gör någonting kommer det att leda till att den tibetanska kulturen dör ut och att det tibetanska folket försvinner . .
( EN ) Jag känner stor sympati för vad ni sade om kulturarv och om den buddhistiska traditionen .
Liksom ni har jag läst Dalai Lamas självbiografi .
Det är en mycket rörande berättelse , inte bara om hans skyldigheter i och gentemot Tibet utan också om hans andliga åskådning .
Kommissionen har , liksom andra , uppmanat till dialog .
Dalai Lama har gjort klart att han önskar en fredlig dialog .
Jag önskar att de kinesiska myndigheterna hade svarat konsekvent och positivt på denna invit från Dalai Lama .
Vid eller omkring tiden för president Clintons besök i Kina gav presidenten i Folkrepubliken Kina intryck av att dialog stod på dagordningen .
Det skulle vara mycket välgörande , inte bara för Tibet och för alla de som tror på fred och stabilitet i Asien , utan det skulle också verkligen vara till heder för Folkrepubliken Kinas regering om den skulle svara på dessa försök att inleda en dialog .
Fråga nr 31 från ( H-0795 / 99 ) : Angående : Stadgan om god förvaltning inom EU som avvisats av kommissionen Enligt uppgifter i pressen har kommissionen avvisat det förslag om medborgarnas rätt till god förvaltning inom EU , vilket framlagts av den europeiska ombudsmannen Jacob Söderman .
Kommissionen har själv godkänt tanken på en stadga för god förvaltning men kom nu att avvisa det detaljerade förslaget och framlade i stället en rad kompletterande föreskrifter om bättre service .
Stämmer de ovannämnda uppgifterna ?
Vad finns det för orsak till att kommissionen handlat som den gjort och hur vill kommissionen förklara den skillnad mellan ord och handling som på det här viset uppstått på tal om förnyandet av EU : s förvaltning ?
Tycker kommissionen att det inträffade stämmer överens med det fempunktsprogram som Europaparlamentet och kommissionen kom överens om i september och är kommissionen beredd att framlägga ett detaljerat förslag till en stadga för god förvaltning i sådan form att också parlamentet har en möjlighet att ta ställning till det ?
Jag överlämnar ordet till Patten , som företrädare för kommissionen . .
( EN ) Den tidningsartikel som ni hänvisar till tycks mig vilseledande och felaktig .
I november 1999 antog kommissionen vid förstabehandling en uppförandekod för tjänstemännen som skulle införlivas med arbetsordningen .
För närvarande rådgör kommissionen med sina tjänstemannarepresentanter om detta dokument , och denna process kommer att slutföras under de närmaste veckorna .
Kommissionen kommer då att anta koden vid andrabehandling .
Man bör notera att den nya kommissionen på eget initiativ omedelbart följde upp den europeiske ombudsmannens beslut från 28 juli 1999 i hans utredning om koden .
Kommissionen skulle speciellt vilja betona att vi när vi upprättade denna kod har anammat alla ombudsmannens förslag till rekommendationer .
Koden kommer att bli ett dokument som uteslutande handlar om kommissionens tjänstemäns förhållande till allmänheten .
Den kommer att antas genom ett juridiskt bindande beslut i kommissionen som kommer att offentliggöras i Europeiska gemenskapernas officiella tidning .
Dokumentet har sammanställts med full hänsyn till de bestämmelser som finns i det förslag som den europeiske ombudsmannens kontor har upprättat .
Enligt bestämmelser i fördragen om detta är det kommissionen själv som ansvarar för att fastställa sin arbetsordning .
Det är emellertid självklart att kommissionen håller fast vid principen om regelbunden politisk dialog med Europaparlamentet om alla aspekter av administrativa reformer .
Herr talman !
Jag vill tacka kommissionären .
Jag frågar ändå , när är det meningen att denna stadga äntligen skall träda i kraft ?
Med tanke på att den har hållit på att utarbetas ända sedan 1997 . .
( EN ) Tidningsartiklarna var vilseledande .
Jag tror inte att det finns någon skillnad mellan oss och ombudsmannen .
Det finns en fråga om den rättsliga grunden och där har vi inhämtat råd och jag tror att vi har väl på fötterna där .
Jag vill upprepa att ledamöter som liksom den ledamot som ställde frågan är speciellt intresserade av denna fråga säkert vill föra en dialog om den .
Det är ytterst viktigt och jag förstår er oro .
Jag vill tacka kommissionen för det som jag uppfattar som ett mycket positivt svar .
För säkerhets skull skulle jag vilja ha en bekräftelse på att det verkligen är så , att det inte finns någon del av Jacob Södermans förslag , vad gäller kommissionen och den goda förvaltningen , som kommissionen tycker är oacceptabel .
Är det korrekt att alla delar av förslaget kommer att godtas till sitt innehåll ? .
( EN ) Låt mig läsa vad det står i mitt sammandrag - och eftersom det står där måste det vara sant !
" Jag skulle återigen vilja betona att kommissionen har godtagit alla ombudsmannens rekommendationer i hans förslag till rekommendationer från juli 1999 " .
Båda dokumenten , det vill säga kommissionens dokument och ombudsmannens förslag , täcker i stort sett samma saker .
Den enda substantiella fråga som har uppstått är den rättsliga grunden .
Jag kan gå in på den i detalj om ni vill men det finns inget tvivel om att vi är ense med ombudsmannen i denna viktiga fråga .
Vi tar gärna med Pattens kommentarer i vår litteraturförteckning , som ett komplement till ledamöternas favoritlektyr .
Eftersom frågeställaren är frånvarande , bortfaller fråga nr 32 .
Jag ber Vitorino om ursäkt för parlamentets ohövliga agerande , vilket jag beklagar .
Enligt arbetsordningen har parlamentet ingen skyldighet att svara .
Jag önskar er en fortsatt bra dag .
Andra delen Frågor till Nielson som har ersatts av Patten Frågorna 33 och 34 i andra delen av frågor till kommissionen är riktade till Nielson .
Nielson kan inte närvara här i dag , eftersom han befinner sig i Sydafrika .
Jag kan meddela att kommissionens vice ordförande Loyola de Palacio har skickat ett brev där hon förklarar detta och meddelar att Patten kommer att vara den som besvarar dessa frågor .
Fråga nr 33 från ( H-0829 / 99 ) : Angående : Mainstreaming i EU-biståndet Ministerrådet utarbetade redan 1995 riktlinjer för integrering av ett jämställdhetstänkande ( mainstreaming ) i hela EU : s biståndspolitik .
Riktlinjerna kräver att all personal som arbetar med utvecklingsfrågor skall få kontinuerlig fortbildning i " gender mainstreaming " , men under de senaste åren har bara ett 50-tal personer utbildats och fortfarande finns ingen obligatorisk jämställdhetsutbildning på generaldirektoratet för bistånd .
Att låta ett jämställdhetstänkande genomsyra den totala verksamheten ( mainstreaming ) innebär att hänsynen till jämställdhet mellan kvinnor och män ingår som en självklar del i alla former av utvecklingspolicy , strategier och insatser .
För att möjliggöra detta måste rådets riktlinjer om mainstreaming tillämpas i sin helhet .
Nuvarande personal måste få obligatorisk utbildning i jämställdhetsfrågor och 1-2 dagars utbildning i jämställdhetsfrågor bör ingå som en nödvändig del i generaldirektoratet för bistånds obligatoriska introduktionskurser för nyanställda .
Är kommissionen beredd att vidta dessa åtgärder ? .
( EN ) Får jag först av allt betona hur ledsen min kollega Nielson var att han inte kunde vara här , men ni som bryr er om dessa utvecklingsfrågor vet säkert hur viktigt hans uppdrag är , att försöka se till att vårt avtal med Sydafrika överlever .
Kommissionen är beredd att titta på möjligheterna att göra en genomgång av jämställdhets- och utvecklingsfrågor till en del av de så kallade introduktionskurserna för ny personal , någonting som redan har förekommit , fast inte regelbundet får jag erkänna .
Utbildning av personal som flyttar till delegationerna i de olika regionerna är en annan inkörsport .
Utbildningen skulle då genomföras automatiskt utan att vara obligatorisk .
Vi siktar också på att lägga in utbildning i dessa frågor i den grundkurs i projektadministration våra tjänstemän genomgår .
Vi vill att detta slags utbildning så långt som möjligt skall vara automatiskt inbyggd i programmen från början i stället för att man skall hantera den separat senare .
Min personliga inställning som före detta utvecklingsminister är att dessa frågor själva borde integreras och tacklas som en del av utbildningen , inte göras till något slags frivilligt tillval .
Strävan efter jämställdhet skall på alla nivåer genomsyra arbetet vid Generaldirektoratet för bistånd .
Den skall inte tillföras som " något vid sidan om " .
Detta måste naturligtvis leda till en omformulering av utvecklingsmål och strategier samt en omvandling av institutioner och processer , så att såväl kvinnors som mäns prioriteringar och behov avspeglas på ett bättre sätt .
Vidare måste åtgärder mot könsgrundade skillnader vidtas .
Jämställdhet måste genomsyra inte bara projekt och program , utan också alla övergripande mål , handlingsplaner och strategier .
Det ser ut som om vi är överens om detta .
Men ansvaret för att vederbörlig uppmärksamhet ägnas jämställdhet ligger hos avdelnings- och enhetschefer .
Om inte cheferna besitter den professionella kompetens som krävs , så sker ingenting - gender mainstreaming bortprioriteras .
Ytterst få i ledningen av Generaldirektoratet för bistånd , dvs. enhetschefer och ännu högre chefer , har deltagit i de genderkurser som har anordnats .
Endast en chef har deltagit i genderutbildningen en halv dag .
Detta är naturligtvis oacceptabelt .
Vad är kommissionen beredd att göra för att se till att enhetschefer och chefer på ännu högre nivå genomgår nödvändig genderutbildning ?
Det har hänt att gender har ingått i den obligatoriska introduktionskursen för nyanställda , men då bara en till två timmar per kurs .
Detta begränsade utbildningsmoment har dock strukits från alla introduktionskurser som har ägt rum under senare tid .
Som jag i min fråga påpekar , krävs det inte att en till två timmar , utan att en till två dagar ägnas åt ämnet .
Min fråga är : Är kommissionen verkligen beredd att fullfölja de antagna riktlinjerna för gender mainstreaming på Generaldirektoratet för bistånd ? .
( EN ) Jag tar verkligen frågan om integrering av ett jämställdhetsperspektiv på allvar , och det gör min kollega kommissionär Nielson också .
Jag skall inte tjata om böcker , men jag har just läst en bok av David Landis Barnhill om vad det är som gör att vissa länder blomstrar och andra inte , och det är intressant att se den betydelse han fäster vid jämställdhetsfrågor för ekonomisk framgång och politisk stabilitet i olika samhällen under årtusendena .
För det andra anser jag att även om den utbildning vi talar om inte bör vara obligatorisk - när allt kommer omkring finns ingen obligatorisk utbildning om någonting hos kommissionen - bör den vara väsentlig .
Och eftersom den bör vara väsentlig skulle man hoppas att alla skulle se till att de hade tillräcklig jämställdhetsutbildning .
Det gäller alla , på alla nivåer .
Det är inte någonting som högre tjänstemän skall bedöma som lämpligt för sina underställda , men tro att de själva är för vuxna eller för högt uppsatta för att genomgå .
För det tredje är ett av de bästa sätten att angripa denna fråga att integrera jämställdheten som en viktig och gränsöverskridande fråga i de mest populära kurserna för utvecklingstjänstemän och framför allt kanske i kursen om projektadministration som är nyckeln till god administration av projekt på fältet .
Så jag håller till stor del med om det ni sade .
Jag hoppas att det angreppssätt vi har anammat visar på både ett praktiskt sinnelag och vikten av att detta får den uppmärksamhet det förtjänar .
Fråga nr 34 från ( H-0831 / 99 ) : Angående : Hjälp åt Centralasien Vilket utvecklingsbistånd och humanitärt bistånd tillhandahåller kommissionen åt staterna i Centralasien , och hur bedömer kommissionen att effekten av detta bistånd är ?
Frågor riktade till Diamantopoulou .
( EN ) Sedan 1991 ger gemenskapen ett betydande ekonomiskt stöd till de nya oberoende staterna och däribland länderna i Centralasien .
Större delen av Europeiska unionens stöd har tillhandahållits inom ramen för Tacis-programmet .
1998 och 1999 erhöll Kirgizistan , Kazakstan , Uzbekistan och Turkmenistan tekniskt bistånd på 75 miljoner euro .
Detta bistånd har gagnat alla områden , särskilt jordbruket , infrastrukturutvecklingen , privatekonomin och stärkandet av institutionerna .
Tadzjikistan har av säkerhetsskäl inte kunnat dra nytta av Tacis fullt ut , men ett återuppbyggnadsprogram på 7,2 miljoner euro har funnits på plats under 1998 och 1999 .
Förutom de nationella programmen har Europeiska unionen stött viktig regional verksamhet inom energi- , transport- och miljösektorerna .
Livsmedelssäkerhetsprogram i Centralasien inleddes 1996 efter att Europeiska unionen under två år levererat livsmedelsstöd in natura .
Dessa program har gagnat Kirgizistan och i mer begränsad omfattning Tadzjikistan .
Avsatta medel för de icke-statliga organisationernas program i Tadzjikistan uppgick till 7,42 miljoner euro 1998 och 1999 .
Under samma period fick Kirgizistan 17 miljoner euro .
Sedan 1993 har kommissionens Europeiska gemenskapernas kontor för humanitärt bistånd , ECHO , aktivt stött de mest utsatta grupperna och sektorerna i Tadzjikistan och Kirgizistan .
För 1998 och 1999 avsattes 3,8 miljoner euro till Kirgizistan och Tadzjikistan erhöll över 35 miljoner euro , huvudsakligen för livsmedel , läkemedel , vatten och hygien .
Det har framgått av regelbundet återkommande utvärderingar och lägesbedömningar att Europeiska unionens stöd bidrar till dessa länders stabilitet och därmed till den pågående fredsprocessen .
Herr talman , herr kommissionär !
Centralasien och Kaspiska havet hotar ju att bli 2000-talets Balkan .
Därför hänger det mycket på en stabilisering av just de stora staterna Turkmenistan och Uzbekistan .
Jag vill därför fråga er , och detta ligger ju inom ert eget ansvarsområde , hur förhandlingarna beträffande partnerskapsavtalet med dessa båda länder går , alltså de politiska förbindelserna .
Det är ju direkt ert område ; min andra fråga gäller kollegan Nielsens område : hur går det ekologiska samarbetet , i synnerhet beträffande vattnet och problematiken med monokulturerna av bomull , som leder till stor uttorkning . .
( EN ) Under toppmötet i Istanbul för några veckor sedan hade vi tillfälle att träffa och föra diskussioner med några av de Centralasiatiska republikerna .
Jag är mycket mån om att vi stärker våra relationer med dem .
Om ni vill kan jag skicka er en detaljerad sammanställning av exakt var vi befinner oss i förhandlingarna om partnerskap och samarbetsavtal med var och en av de Centralasiatiska republikerna .
Alla hoppas naturligtvis att denna förutsägelse om vad som kan hända i framtiden är för pessimistisk .
Men jag tvivlar inte alls på att ni har rätt när ni betonar Centralasiens strategiska betydelse .
Jag har tidigare hört er tala om Kaukasus också .
Ni har helt rätt i att en union som talar om att förhindra konflikter borde titta på vad den kan göra i dessa speciella områden för att tillse att den typ av konflikt inte uppstår som den på Balkan som har orsakat så mycket förödelse och som har kostat oss en hel del mer än vi kanske skulle ha gjort av med annars , om vi hade vidtagit fler förebyggande åtgärder , om dessa hade varit möjliga .
Så era kommentarer om dessa regioners strategiska betydelse är ytterst välfunna .
Vi bidrar till program i regionen som har viss miljöpåverkan .
Våra livsmedelsprogram hänger direkt samman med strukturella jordbruksreformer liksom med lindrande av fattigdom .
Dessa program syftar i sig till att säkerställa att jordbruket får en sundare bas i dessa samhällen och inte bara går ut på att våldta jorden .
Det finns en ekologisk aspekt som vi bör fortsätta att prioritera .
Lägg märke till att den ledamot som ställde frågan applåderade kommissionärens svar .
Det sker inte så ofta .
Och dessutom har kommissionären i det här fallet inte nämnt litteraturförteckningen .
Tack så mycket , herr Patten , för era inlägg i dag .
Fråga nr 35 från ( H-0778 / 99 ) : Angående : Greklands åtgärdsplan för sysselsättningen Enligt vad som framkommit vid utvärderingen av åtgärdsplanerna för sysselsättning har kommissionens kritik huvudsakligen riktats mot Grekland och Italien för att dessa inte på vederbörligt sätt genomfört sysselsättningspolitiken och stödåtgärderna för sysselsättningen .
I rapporten konstateras det att varken Grekland eller Italien ännu nått målen för förbättrad anställbarhet och att det är tvivel underkastat om den politik som avses genomföras kommer att göra det möjligt att följa riktlinjerna för hur långtidsarbetslösheten skall förebyggas eller hanteras .
I rapporten ingår också en kommentar om att Grekland inte planerat några åtgärder på medellång eller lång sikt för att sänka arbetsgivarens skatter och försäkringsavgifter i samband med anställande och att det dessutom inte föreligger några exakta siffror över sysselsättningen .
Kan kommissionen upplysa om Greklands regering ingått några särskilda åtaganden för hur problemet med ungdoms- och långtidsarbetslöshet kunde angripas och vilka dessa åtaganden i så fall är ?
Har regeringen lagstiftat om och infört något system för hur växlingarna i sysselsättning skall kunna fastställas , registreras och övervakas eller handlar merparten åtgärder fortfarande bara om att räkna dem som är utan arbete ?
Som svar på Papayannakis fråga kan jag säga att det i åtgärdspaketet för sysselsättning 1999 framförde kommissionen vissa förslag och rekommendationer till Grekland i syfte att effektivisera sysselsättningsåtgärderna .
Den viktigaste punkten var att man måste anstränga sig för att reformera den offentliga förvaltningen , där det finns problem .
Man måste förbättra systemet för statistisk uppföljning och vidta förebyggande politiska åtgärder i enlighet med riktlinjerna 1 och 2 i sysselsättningspaketet .
Jag måste tala om att den grekiska regeringen , inom ramen för sin arbetslöshetspolitik , har två konkreta program för 1999 : " ja till yrkeslivet " och " tillbaka till arbetet " .
Jag har ännu inte fått veta det slutliga resultatet av dessa program , så att jag kan se om de kvantitativa målen har uppnåtts .
Den grekiska regeringen är i dag medveten om problemet med att man inte kan registrera flödet av arbetskraft till och från sysselsättning och har därför åtagit sig , för det första , att omorganisera landets arbetsmarknadsmyndigheter , för det andra , att skapa effektiva centra för främjande av sysselsättning - detta program har redan inletts men har ännu inte avslutats - för det tredje , att införa ett lämpligt system för elektronisk registrering av sysselsättningen för att kunna följa upp alla dessa praktiska åtgärder .
I det nya programmet för perioden 2000-2006 , som finansieras av Europeiska socialfonden , bör man , även med kommissionens stöd , utnyttja alla nödvändiga resurser och politiska åtgärder för att förverkliga de mål jag tidigare nämnde .
Kommissionen kommer att noga följa hur den grekiska regeringen fullföljer sina åtaganden .
Jag tackar kommissionsledamoten för hennes svar .
Men , fru kommissionär , vi befinner oss i följande situation .
I fråga om arbetslöshetens omfattning ligger vi på andra plats i Europa , dvs .
11,3 procent - vilket vi inte gjorde tidigare - , vi har den största ökningen av arbetslösheten , vi lägger ut minst pengar på de arbetslösa , dvs. mindre än 1 procent av BNP , medan andra länder spenderar 3-4 procent ( t.ex.
Frankrike , Belgien och Tyskland ) , och det är inte klart hur man har använt de pengar som Europeiska socialfonden betalat ut , bl.a. för att bekämpa arbetslösheten .
Ni säger att kommissionen har lämnat vissa rekommendationer .
Jag gläder mig över detta och hoppas att man följer rekommendationerna .
Men jag har väldigt länge burit på en fråga : hur har det gått med de tidigare politiska åtgärderna ?
Är det någon som fått ett arbete ?
Hur många har fått arbete ?
I fjol och i förfjol , om ni inte kan säga hur det är i år .
Hur har det gått med yrkesutbildningen ?
Dessa så omtalade utbildningscentra , är de till för att ge arbete åt dem som utbildar eller åt dem som utbildas ?
Har vi några siffror ?
Har vi således någon möjlighet att kontrollera hur den grekiska regeringen sköter denna politik ?
Herr Papayannakis !
Vad jag skulle kunna svara är att vad den grekiska regeringen verkligen bör satsa på är den elektroniska statistiska registreringen av befintliga strukturer , så att de pågående programmen kan ge de kvantitativa resultat som ni talar om , men också för att möjliggöra en uppföljning som ger underlag för den politik som bör föras .
Grekland har uppvisat en ökad sysselsättningsgrad och - efter vad jag kan se här - också en ökad produktivitet .
Det kommissionen kan påverka är de konkreta riktlinjerna .
Som ni vet , är det 22 riktlinjer som varje land bedöms efter .
De gäller tillgång till yrkesutbildning och de speciella åtgärderna för långtidsarbetslösa .
I fråga om alla dessa riktlinjer kommer kommissionen att försöka få fram kvantifierbara data och konkreta uppgifter om förverkligandet av gemenskapens riktlinjer för perioden 2000-2006 .
Fråga nr 36 från ( H-0782 / 99 ) : Angående : Det danska systemet för förtidspension Har kommissionen godkänt det danska systemet för förtidspension i sin helhet ?
Råder det eventuell oenighet mellan Danmark och kommissionen på andra socialpolitiska områden ?
Det danska pensionssystemet , Eftarløn , innebär att pension endast kan utgå till dem som är bosatta i Danmark och till dem som uppfyller kravet på att ha arbetat en viss tid i detta land .
Det finns arbetstagare som framfört klagomål till Europeiska kommissionen för att de inte har rätt till pension .
De danska myndigheterna anser inte att gemenskapslagstiftningen tvingar dem att betala ut denna ersättning till förtidspensionerade arbetstagare , när dessa inte uppfyller villkoren enligt dansk lag .
Det bör noteras att gällande förordning om socialförsäkringssystem för närvarande inte omfattar några bestämmelser om förtidspensionering , och kommissionen har föreslagit vissa förändringar i förordningen , vilka emellertid ännu inte har avgjorts av rådet .
EG-domstolen har hittills ännu inte tagit ställning till Eftarløn , men man skulle på goda grunder kunna hävda att bosättningsvillkoren inte är förenliga med de allmänna kraven på förbud mot diskriminering på grund av medborgarskap .
Europeiska kommissionens tjänsteenheter har inlett ett förfarande med möten och överläggningar med den danska regeringen för att kunna nå fram till en gemensam lösning .
Det senaste mötet i denna fråga hölls i november 1999 , och vi avvaktar slutliga förslag från kommissionens tjänsteenheter om huruvida det kan bli aktuellt med ett ingripande mot Danmark .
Jag lade märke till att kommissionsledamoten inte gav något direkt svar på frågan om det danska förtidspensioneringssystemet i sin helhet är godkänt av kommissionen , men det framgick ju indirekt att svaret var nekande .
Jag vill be kommissionsledamoten att uttryckligen bekräfta att systemet inte är godkänt av kommissionen .
Kommissionen gjorde ju mer än bara antydde att man starkt överväger att ta upp hela frågan om det danska förtidspensioneringssystemet i domstolen i Luxemburg , just med den utgångspunkt att det här föreligger en faktisk diskriminering i förhållande till icke-danska arbetstagare som inte kan uppfylla villkoren till följd av att de inte arbetat under den tidsperiod som krävs enligt det danska systemet .
Jag vill fråga kommissionären om hon kan ange några ungefärliga tidsperioder i detta sammanhang , eftersom det är ett problem som måste få ett avgörande i den danska socialpolitiska debatten .
Jag skulle alltså vara tacksam om kommissionären skulle kunna utveckla denna fråga .
Herr parlamentsledamot !
Vad jag skulle vilja framhålla är att det såväl i Danmark som i många andra länder finns problem i fråga om tolkningen av direktiven , när de skall införlivas med respektive lands lagstiftning .
Detta är ett sådant fall. och det pågår en diskussion mellan den danska regeringen och kommissionen , för att frågan skall kunna lösas på bästa sätt , till gagn för de arbetstagare som uppfyller villkoren och som , enligt gällande lagstiftning , har denna rätt till pension .
För att bara helt kort knyta an till den sista punkten .
Jag uppmanar kommissionen att göra det helt klart att kommissionens invändningar , för vad de är värda , inte på något sätt skulle inkräkta på danska medborgares rätt att dra nytta av denna plan utan att kommissionen bara är angelägen , vilket den har rätt att vara enligt gemenskapens lagar , om att säkerställa att planen gäller alla gemenskapsmedborgare som uppfyller villkoren .
Jag anser att svaret är kort och tydligt .
Det är naturligtvis så som ni sade .
Det kommer inte att bli något problem med de danska medborgarna , och det är inte där problemet ligger .
Problemet gäller danska eller andra medborgare , som är bosatta utanför Danmark .
Fråga nr 37 från ( H-0791 / 99 ) : Angående : Arbetstidsdirektivet Sjukhusläkare , som inte är konsulterande , omfattas inte av arbetstidsdirektivet från 1993 och inte heller av förslaget till ändring av rådets direktiv ( KOM ( 98 ) 0662 - C4-0715 / 98-98 / 0318 ( SYN ) ) .
Vilka åtgärder föreslår kommissionen för att säkerställa att skyddsnivån för dessa läkare är jämförbar med den som fastställs i direktivet från 1993 ?
Fråga nr 38 från ( H-0805 / 99 ) : Angående : Åtgärder för att öka jämställdheten mellan könen En av de arbetsgrupper av kommissionsledamöter som har aviserats av ordförande Prodi har som mål att främja åtgärder för ökad jämställdhet mellan könen ( införlivande av jämställdhetsaspekten , så kallad mainstreaming ) .
Vilka kommissionsledamöter ingår i denna grupp ?
Hur många gånger har de träffats hittills ?
Vilka konkreta åtgärder har diskuterats ?
Frågan innehåller flera delfrågor .
Den gäller kommissionens särskilda kommitté som sysslar med jämställdhetsfrågor .
De kommissionsledamöter som medverkar är ordföranden Prodi , vice ordföranden Kinnock , Reading och jag själv .
Kommitténs sammanträden är öppna , och det första sammanträdet hölls den 11 januari 2000 .
Vi diskuterade tre allvarliga frågor : den första gällde det femte kvinnoprogrammet , som vi efter min föredragning hade en första diskussion om , den andra gällde Busquins rapport om undersökningen av kvinnors deltagande i forskning och vetenskap , och den tredje gällde Kinnock , som informerade kommissionen om ansträngningarna att ta hänsyn till jämställdhetsaspekten i det omfattande reformarbete som i dag pågår inom gemenskapen .
Tack för ert svar , fru kommissionär , men jag måste beklaga att det dröjde så länge innan arbetsgruppen kom samman , med tanke på hur viktig den här frågan är , och vi litade på att den här kommissionen redan från starten skulle börja eftersträva en större jämlikhet mellan kvinnor och män .
Jag hoppas att det kommer att ske en förändring och att sammankomsterna blir täta , för det finns många frågor som kommissionen måste ta itu med , så att de åtgärder som leder till en större jämlikhet mellan kvinnor och män påskyndas och leder till goda resultat så snart som möjligt .
Fru ledamot , här rör det sig om en uppmaning och inte om en fråga .
Men om fru kommissionären vill ge någon förklaring eller visa sin goda vilja ...
Låt mig bara få säga en sak till : jag håller med om att kommissionen borde ha sammanträtt tidigare , men förseningen kompenseras av innehållet i sammanträdet , för vi fattade genast viktiga beslut .
Fråga nr 39 från ( H-0807 / 99 ) : Angående : Gemenskapsinitiativet Equal Den 13 oktober 1999 antog kommissionen gemenskapsinitiativet Equal som syftar till att främja gränsöverskridande samarbete och till att finna och utveckla nya sätt att bekämpa diskriminering och ojämlikhet som på arbetsmarknaden .
Initiativet är främst inriktat på asylsökande .
Inom ramen för detta initiativ skall varje medlemsstat lägga fram förslag i form av ett gemenskapsinitiativ som omfattar den egna staten .
Vilka kriterier kommer kommissionen att grunda sig på för att godkänna eller avslå medlemsstaternas föreslagna program ?
Vilket gemenskapsorgan skall kontrollera finansieringen av den verkställande kommittén och uppföljningskommittén , och att programmet genomförs på ett riktigt och oklanderligt sätt ?
Anslagen från Europeiska socialfonden kommer för perioden 2000-2006 totalt att uppgå till 2,487 miljarder euro .
Hur mycket kommer Grekland själv att bidra med tanke på att gemenskapsinitiativet Equal är ett initiativ som förutsätter samfinansiering från medlemsstaternas sida ?
Initiativet Equqal är inte begränsat till vissa grupper av människor .
Det gäller hur man skall motverka diskriminering på arbetsplatserna .
Beslutet om detta initiativ fattades i Berlin , och då beslutade man att det även skall omfatta de yrkesarbetande bland dem som söker asyl .
Jag vill framhålla detta som ett viktigt inslag i detta direktiv .
I varje medlemsstat måste gemenskapsinitiativets program överensstämma med de stadgar som gäller Europeiska socialfonden , dvs .
Equqal följer socialfondens stadgar .
Det har presenterats för parlamentet , och vi väntar på parlamentets yttrande i nästa månad .
Jag måste betona att initiativet Equal svarar mot nationella behov och nationell planering i enlighet med den överenskomna europeiska strategin .
Det är i första hand de nationella regeringarna som har ansvaret för att inrätta de gemensamma organen och lägga fram förslag och utse dem som skall genomföra programmen , men det är också i första hand de nationella regeringarna som skall ansvara för kontrollen .
Inom Europeiska kommissionen finns Generaldirektoratet för sysselsättning , som ansvarar för genomförandet , och budgetkontrollen utövas av Generaldirektoratet för budgetkontroll , av Europeiska byrån för bedrägeribekämpning och av Europeiska revisionsrätten .
Slutligen har vi frågan om vilken summa som har betalats ut .
Grekland har fått 98 miljoner ecu med krav på 80 procents medfinansiering .
För öregionerna och framför allt för de mest avlägset belägna grekiska öarna uppgår initiativets andel till 85 procent och medfinansieringen uppgår till 15 procent .
Herr talman !
Jag anser att riktlinjerna för gemenskapsinitiativet Equal , och speciellt de fyra åtgärder som beskrivs i det , leder till ett mycket komplicerat , byråkratiskt , men egendomligt nog också svåröverskådligt system .
Man frågar sig t.ex. på vilket sätt ett utvecklingssamarbete skall bevisa att det är representativt och präglas av samarbetsanda , såsom krävs av åtgärd 2 i artikel 33 i direktiven .
Kravet på mellanstatligt samarbete och de komplicerade kraven på planering och genomförande av ett utvecklingssamarbete leder ofrånkomligt tanken till stora system , som ensamma kan uppfylla dessa krav .
Detta strider emellertid mot de allmänna målens uttalade önskemål om decentraliserade handlingsplaner , helst på den lokala självstyrelsens eller jordbruksområdenas nivå .
När det gäller de mest utsatta grupperna , såsom asylsökande , invandrare och andra , innebär det att deras medverkan är omöjlig eller bara symbolisk .
Om man tänker på att den totala summan är ganska liten - 2,8 miljarder euro för så ambitiösa mål i 15 stater - är jag rädd att det enda vi till sist kommer att kunna bevisa är att arbetslösheten är av ondo .
Först skulle jag vilja säga att det skulle vara till stor hjälp för mig , när vi nu behandlar frågan i parlamentet , om ni ville framföra konkreta förslag , som jag kan ta ställning till .
För det andra måste jag säga att initiativet Equal varken avser eller kan minska arbetslösheten eller stödja sysselsättningsfrämjande åtgärder .
För detta ändamål finns den europeiska sysselsättningsstrategin och Europeiska socialfonden , som förfogar över mycket stora summor och utomordentligt stora resurser , i synnerhet för länder som Grekland .
Initiativet Equal har en konkret uppgift .
Att hjälpa till med att få fram statistiskt material , att genomföra undersökningar och inrätta organ som skall kunna stödja de grupper inom befolkningen som drabbats av diskriminering .
Vad vi eftersträvar är alltså samarbete mellan lokala grupper , organ för lokal självstyrelse , mellan länder , så att ett erfarenhetsutbyte kommer till stånd .
Vi vill alltså framför allt att länderna skall utbyta erfarenheter med varandra .
Det är dessa tankar som ligger till grund för initiativet och som också avspeglas i dess budget .
Vårt mål är att samarbetet i största möjliga utsträckning skall omfatta utvecklingsprogram , privata organisationer , lokala myndigheter , för att komma så nära medborgarna som möjligt .
Fråga nr 40 från ( H-0808 / 99 ) : Angående : Artikel 13 i EU-fördraget och sysselsättning Det förslag till kommissionens direktiv som fastställer en allmän ram för likabehandling inom ramen för anställning och sysselsättning , beviljar undantag för religiösa organisationer ( artikel 4.2 ) .
Kan kommissionen informera parlamentet om vilka situationer och grupper inom ramen för artikel 13 ( EU-fördraget ) som kan påverkas av ett sådant undantag ?
För en månad sedan lade kommissionen fram ett förslag i frågan om lika behandling i arbetslivet , i överensstämmelse med fördragets uppdrag att genomföra artikel 13 .
Förbud mot diskriminering är ledstjärnan i vårt paket med direktiv och program .
Men efter förslag från kommissionen och efter ungefär två års överläggningar med arbetsmarknadens parter , med medlemsstaterna , med Europaparlamentet , finns det vissa undantag .
Och dessa undantag gäller de yrken som måste utövas av personer med en specialiserad yrkesutbildning .
Och jag kan ge ett mycket konkret exempel för att förtydliga .
I en religiös skola är det rimligt att man begär och beviljas undantag , med innebörden att den lärare som tjänstgör vid den aktuella skolan skall omfatta samma konfession som skolan .
Undantagen är alltså av detta slag .
Det rör sig inte om generella undantag , utan dessa skillnader i fråga om behandling i enlighet med de olika medlemsstaternas specialbestämmelser är berättigade endast när det gäller denna specialiserade yrkesutbildning .
Detta är en snedvriden tolkning av hur man stoppar diskriminering .
Till exempel skulle det vara helt i sin ordning om religiösa skolor sade till en katolik : vi vill inte anställa dig för du är homosexuell .
Det vi har här från kommissionen är en förstärkning av en förtryckande hierarki .
Det vi borde göra är ju , och jag hoppas ni instämmer herr kommissionär , att anställa människor på grundval av deras kompetens och inte bevara ett sådant bigotteri och en sådan fördomsfullhet , oavsett hur starkt övertygad man än är. kommissionen .
( EL ) Jag vill betona att detta undantag inte innebär att man kan vägra en person anställning av vilket skäl som helst .
Av det skäl ni nämnde , på grund av sexuell läggning , etnisk diskriminering eller vad det vara månde .
Undantaget ger en möjlighet till urval endast i de fall då det krävs speciell kompetens , som har ett direkt samband med verksamheten .
Det är alltså fråga om positiv diskriminering .
I det exempel ni nämnde , i den katolska skolan , är det logiskt att läraren skall vara katolik .
Det är bara undantag av detta slag som kan accepteras .
Fråga nr 41 från ( H-0813 / 99 ) : Angående : Främjande av sysselsättning för kvinnor i starkt missgynnade regioner Kvinnor som lever i starkt missgynnade regioner har ofta enorma svårigheter att få arbete .
De har i många fall inte något minimikapital och i deras miljö saknas företagaranda , kooperativa traditioner och utbildningsmöjligheter .
De är dessutom bosatta i landsbygdsområden där 80 procent av befolkningen befinner sig nära fattigdomsgränsen .
Vilka åtgärder planeras för att hjälpa dessa kvinnor att överbrygga hinder som hänger samman med deras sociala bakgrund ?
Har kommissionen för avsikt att lägga fram en politik som säkerställer en miniminivå , för att på ett korrekt sätt återspegla de extrema förhållanden som dessa kvinnor faktiskt lever under , eller kommer deras svåra situation att återigen förbigås i den nya sysselsättningspolitiken ?
För de eftersatta områdena i Europa finns ju sammanhållningspolitiken , och för att genomföra denna politik finns samarbetet och de gemensamma insatserna av både strukturfonderna och Europeiska socialfonden och jordbruksfonden .
Jag vill tala om att de tillgängliga resurserna för problemområdena utgör en tredjedel av den totala budgeten .
Dessa regionalpolitiska insatser som utförs enligt gemensamt överenskomna europeiska riktlinjer i varje medlemsstat - dvs. varje medlemsstat har ansvaret för att genomföra detta program - syftar till att öka antalet arbetstillfällen för både män och kvinnor .
Jag kan tala om att 70 procent av bidragen för perioden 2000-2006 , som uppgår till 195 miljarder euro , kommer att gå till de mest eftersatta regionerna i Europa .
När det nu speciellt gäller kvinnornas möjligheter till förvärvsarbete , vill jag säga , för det första , att socialfonden innehåller en hel pelare med åtgärder som medlemsstaterna måste vidta för att skapa jämställdhet i fråga om arbetstillfällen , dvs. speciella politiska åtgärder som finansieras av socialfonden och gäller kvinnor .
För det andra , i initiativet Leader , som just nu är föremål för granskning , prioriterar man särskilt de utvecklingsstrategier som speciellt syftar till att stödja kvinnor i småföretag inom jordbrukssektorn , inom agroturismen , för att sysselsättningen för kvinnor i jordbruksområdena skall öka .
Tack fru kommissionär .
Ni har gett mig ett välment och precist svar i ordalag som jag uppskattar .
Ändå kan jag försäkra er om att vi med de medel som finns tillgängliga - och som ni nämner - inte kan nå de missgynnade regionerna .
För det är regioner där bristerna tar överhanden , och de bör likställas med sådana regioner där vi arbetar i ett partnerskap , där det i princip råder brist på allting .
Därför undrar jag om ni inte kan undersöka möjligheten att politiken med mikrokrediter , som har gett resultat för partnerskapet , kan tillämpas bland kvinnor i starkt missgynnade regioner , där de har alla odds emot sig .
Jag känner väl till de program ni nämner .
Jag kan försäkra er om att vi med hjälp av dessa inte når dit där behoven är som störst .
Med hjälp av strukturpolitiken - som jag är väl förtrogen med - och med Leader och utvecklingen på landsbygden kan vi inte , vilket behövs , främja sysselsättningen bland kvinnor i de missgynnade regionerna .
Därför ber jag att ni undersöker möjligheten att en politik med mikrokrediter tillämpas .
Kommissionären instämmer och lovat att lägga Izquierdo Rojos anförande på minnet .
Fråga nr 42 från ( H-0817 / 99 ) : Angående : Kommissionens planer beträffande presenterandet av ett nytt socialt handlingsprogram Det är angeläget att kommissionen snarast presenterar ett nytt socialt handlingsprogram vari en konkret plan redovisas , inklusive tidtabell för genomförande för såväl det lagstiftande arbetet inom området för social trygghet som initiativ till ramavtal inom ramen för den sociala dialogen .
Kan kommissionen redogöra för sina konkreta avsikter vad gäller framläggandet av ett nytt socialt handlingsprogram ?
Jag räknar med att det nya programmet för kommissionens socialpolitik under nästa femårsperiod kommer att vara färdigt i slutet av sommaren år 2000 .
För att detta program skall bli färdigt och för att vi skall kunna presentera det , bör vi först slutföra överläggningarna med parlamentet , med arbetsmarknadens parter och med de icke-statliga organisationerna .
Det är en diskussion som börjar nu , men vi bör ta hänsyn till resultaten från Lissabonmötet .
Vid Europeiska rådets möte i Lissabon görs ett nytt försök att ta itu med frågan om den sociala utslagningen , den sociala utslagningens samband med informationssamhället , med den ekonomiska politiken och med reformerna .
Dessa resultat kommer att vara mycket viktiga för den slutliga utformningen av kommissionens sociala program .
Jag har redan tidigare nämnt för Europaparlamentet att ett möte mellan parlamentet och kommissionen kommer att hållas efter Lissabonmötet för att diskutera alla aspekter i fråga om den slutliga utformningen av det sociala programmet för perioden 2000-2006 .
Det är klart att ett kommande socialt handlingsprogram skall ta hänsyn till utvecklingen , t.ex. inom informationsteknologin , och vara ett modernt socialt handlingsprogram i tiden .
Men kan ni också bekräfta det som jag tar upp i min fråga , nämligen att programmet kommer att få en sådan utformning att vi får en konkret tidtabell för de olika typer av lagstiftning på det sociala området , som kommissionen planerar , samt för de initiativ som kommissionen planerar när det gäller den sociala dialogen mellan arbetsmarknadens parter .
Vi har ett behov av att se vilka konkreta alternativ kommissionen kommer att ta upp under den kommande perioden och vilka initiativ till avtal den kommer att ta .
Jag delar helt er uppfattning , för det första , om att man skall ta hänsyn till informationssamhället - det nämnde jag också .
Den sociala utslagningen , kvinnoprogrammet , våra satsningar i fråga om de sociala trygghetssystemen , allt detta måste man nu betrakta ur det nya perspektiv som informationssamhället innebär .
För det andra ; för de initiativ som tas kommer det naturligtvis att finnas en tidsplan för genomförande och systematisk uppföljning .
Det finns en punkt där jag inte kan göra några bindande uttalanden , och det gäller lagstiftningen på socialförsäkringsområdet .
Som ni vet , omfattas denna inte av fördragets artiklar , dvs. fördraget innehåller ingen rättslig grund för socialförsäkringsområdet .
Eftersom frågeställaren är frånvarande bortfaller fråga nr 43 .
Fråga nr 44 från ( H-0819 / 99 ) : Angående : Handikappades möjligheter att ta del av den fria rörligheten inom EU I enlighet med artikel 13 Amsterdamfördraget skall varje EU-medborgare kunna ta del av den fria rörligheten inom unionen .
För personer med olika slags fysiska handikapp , i behov av särskilda transporter och personlig assistans , är dock denna fria rörlighet fortfarande mycket begränsad .
Vilka åtgärder vidtar kommissionen för att underlätta de handikappades möjligheter på detta område ?
Den 26 november 1999 godkände Europeiska kommissionen ett åtgärdspaket för bekämpning av diskriminering .
När det gäller detta paket och personer med funktionshinder , finns det ett direktiv , som går ut på att bekämpa diskriminering , speciellt på arbetsplatserna .
Europeiska kommissionen tror att detta initiativ för bekämpning av diskriminering kommer att bidra till en högre sysselsättningsgrad för personer med funktionshinder och slutligen kommer att underlätta dessa personers fria rörlighet .
Det är naturligtvis särskilt viktigt att personer med funktionshinder får tillgång till kommunikationer , myndigheter och alla slags inrättningar , så att personer med funktionshinder får möjlighet till fri rörlighet .
Europeiska kommissionen har godkänt ett förslag till direktiv om specialbestämmelser för bussar , långfärdsbussar och andra fordon , så att dessa blir tillgängliga även för rörelsehindrade personer , inklusive rullstolsburna .
Dessutom kan jag meddela att rådet den 4 juni 1998 godkände en rekommendation om att införa en typ av alleuropeiskt parkeringskort för personer med funktionshinder , och syftet med rekommendationen är att hjälpa dem att röra sig fritt i alla medlemsländerna med hjälp av ett gemensamt parkeringskort , så att de kan utnyttja alla anordnade parkeringsplatser i Europa .
Jag tackar kommissionären för svaret .
Min fråga rör i första hand handikappades möjligheter att passera gränserna i Europa .
Det är en ganska dyr historia om man skall ta sig från Göteborg till någon plats i övriga Europa på semester eller på studiebesök om man sitter i rullstol och dessutom behöver ha med sig en personlig assistent eller medhjälpare för att klara av situationen .
Jag är tacksam över att kommissionen har antagit en handlingsplan .
Det är ju emellertid en förutsättning att det finns ekonomiska resurser och möjligheter att rent fysiskt komma över gränserna om man har ett funktionshinder .
Det skulle vara intressant att höra om kommissionen också är beredd att avsätta ekonomiska medel för de personer som har funktionshinder , så att också de skall kunna ta sig längre ut i världen än dit rullstolen tar dem .
Jag nämnde kommissionens förslag till direktiv om att de allmänna kommunikationerna måste utformas så att de kan utnyttjas av personer med funktionshinder .
Rådet har inte tagit ställning till förslaget , som är föremål för överläggningar .
Jag anser att ett sådant strategiskt beslut kan fattas på europeisk nivå .
Det är enligt min mening utomordentligt svårt med en specialinriktning för att lösa varje enskild persons transportproblem .
Detta oavsett om det gäller specialprogrammen för utbildning , för ungdomar och kvinnor eller om det måste genomföras genom nationell politik .
Fråga nr 45 från ( H-0006 / 00 ) : Angående : Genomförande av direktiv 96 / 71 / EG om utstationering av arbetstagare Direktivet om utstationering har ännu inte genomförts i Danmark trots att tidsfristen har löpt ut .
Det lagförslag som lagts fram i folketinget innehåller inga bestämmelser som reglerar lönearbetsrättigheter enligt kollektivavtal .
Enligt artikel 3.8 i direktivet skall arbets- och anställningsvillkor vara i överensstämmelse med de " kollektivavtal som har ingåtts av de mest representativa arbetsmarknadsorganisationerna på nationell nivå och som gäller inom hela det nationella territoriet " .
En sådan användning av ett avtal utanför dess individuella område kan emellertid inte åläggas parterna utan stöd i lagen .
Det finns därför två möjliga lösningar : antingen gäller direktivet inte i Danmark eller så innebär direktivet att Danmark måste införa allmängiltiga avtal .
Kan kommissionen bekräfta att direktivet om utstationering inte gäller i Danmark beträffande " kollektivavtal " med " allmän giltighet " ( se artikel 3.1 ) eftersom sådana avtal med allmän giltighet inte existerar i dansk rätt ?
Om inte , hur skall direktivet uppfyllas på denna punkt ?
Europeiska unionens direktiv om utlandsplacering av arbetstagare innebär att samma arbetsvillkor som gäller för mottagarlandet också skall gälla för de utländska arbetstagare som placerats i detta land .
Direktivet innebär att två regelsystem kan tillämpas : antingen mottagarlandets lagstiftning eller de kollektivavtal som tillämpas generellt inom en viss bransch .
Eftersom Danmark inte har ett system som innebär att kollektivavtal upphöjs till allmänt gällande regler , måste man vid tillämpningen av lagstiftningen räkna med att inte bara lagstiftningen om arbetsvillkor utan också de allmänt tillämpliga kollektivavtal som slutits av de mest representativa organisationerna gäller för de utlandsplacerade arbetstagarna .
Enkelt uttryckt kan man alltså säga att Danmark har två alternativ ; antingen att stifta lagar eller också att välja ut ett kollektivavtal och ge det status av lag .
Det förs en diskussion mellan Europeiska kommissionen och Danmark , och vi räknar med att Danmark skall meddela när detta direktiv har införlivats i dess nationella lagstiftning .
Danmarks tidsfrist för att besvara kommissionens frågor löpte ut den 6 december 1999 .
Vi har inte fått något svar .
Vi avvaktar för att se vilka steg som kommer att tas i fortsättningen .
Tack för ett mycket tydligt svar som - om tolkningen stämmer - innebär att direktivet om utstationering medför en skyldighet för danska staten att inrätta ett system med allmänt användbara avtal .
Det är ett mycket tydligt svar , men det är också ett svar - vilket jag måste göra er uppmärksam på - som ställer de danska organisationerna , den danska regeringen och det danska folketinget i en politiskt sett mycket , mycket svår situation , eftersom det är känt att det finns några grundläggande problem i förhållandet mellan den danska modellen som i hög grad bygger på kollektiva avtal , och den kontinentala modellen som förutsätter lagstiftning .
Den oenighet och korrespondens som ni , fru kommissionsledamot , hänvisar till , rör ju först och främst ett annat direktiv , dvs. arbetstidsdirektivet , men nu kan vi alltså se fram emot en ny uppmaningsskrivelse och kommande domstolsförhandlingar som ett resultat av att den danska regeringen inte kommer att , eller uttryckligen har meddelat , att man inte har för avsikt att genomföra lagstiftning och tillämpa allmänt användbara avtal .
För det första ; vi försöker inte ändra systemet vare sig i Danmark eller i något annat land .
Som jag svarade tidigare , finns det alltid problem när det gäller tolkningen av Europeiska kommissionens direktiv , dels därför att de är mycket allmänt hållna , men dels också därför att systemen skiljer sig mycket mellan de olika länderna .
När det gäller er fråga , kan jag säga att det konkreta problemet inte bara gäller Danmark .
Det är inte bara Danmark som har olösta frågor .
Fem länder har införlivat direktivet i sin nationella lagstiftning , och i de övriga pågår diskussioner .
Det har förts diskussioner mellan kommissionen och den danska regeringen men också de andra regeringarna , därför att man måste hitta den bästa metoden för att utlandsplacerade arbetstagare i Danmark skall omfattas av beslut som fattats på europeisk nivå av alla medlemsländerna .
Vi räknar med att både Danmarks och ytterligare nio länders regeringar skall vidta åtgärder i denna riktning .
Tack fru kommissionär för det engagemang ni har visat .
Ni har lyckats uppnå dagens mål : att besvara samtliga frågar .
Vi gratulerar er till detta .
Eftersom tiden för frågestunden med frågor till kommissionen är över , kommer frågorna nr 46 och 68 att besvaras skriftligen .
Jag förklarar härmed frågestunden avslutad .
( Sammanträdet avbröts kl .
19.50 och återupptogs kl .
21.00 . )
 
Ansvarsfrihet 1997 Nästa punkt på föredragningslistan är betänkande ( A5-0004 / 2000 ) av van der Laan för budgetkontrollutskottet om beviljande av ansvarsfrihet för kommissionen och om avslutningen av räkenskaperna för Europeiska gemenskapernas allmänna budget för budgetåret 1997 ( avsnitten I - Parlamentet , II - Rådet , III - Kommissionen , IV - Domstolen , V - Revisionsrätten ) ( SEK ( 1998 ) 520 - C4-0350 / 1998 , SEK ( 1998 ) 522 - C4-0351 / 1998 , SEK ( 1998 ) 519 - C4-0352 / 1999 ) .
Kommissionären är ännu inte här , men jag hoppas och antar att hon kommer om ett par minuter .
Jag vill föreslå att vi börjar trots detta , och hoppas att kommissionären , om hon fortfarande är kvar på sitt kontor , kan lyssna till talet , i synnerhet föredragandens tal .
Herr talman !
Fru Schreyer har säkerligen ett mycket gott skäl för att inte vara här , för annars skulle hennes frånvaro vara oförlåtlig .
Jag skulle vilja börja med att tacka mina kolleger för deras medverkan till detta betänkande .
Det skulle inte ha varit vad det är i dag utan denna samarbetsanda .
Herr talman !
I början av förra året sköts beviljandet av ansvarsfriheten för 1997 upp , eftersom parlamentet omöjligen kunde bevilja ansvarsfrihet åt en avgående kommission som inte skulle kunna åta sig förpliktelser för framtiden .
I sin resolution hävdade parlamentet att ansvarsfrihet skulle kunna beviljas först efter det att vi fått seriösa , långtgående reformförslag från den nya Europeiska kommissionen .
Detta betänkande läggs nu fram vid en avgörande tidpunkt , omedelbart före Kinnocks reformer .
Det är en utmärkt chans för parlamentet att sätta en långtgående reformstämpel på dessa planer .
Redan under förarbetet har det visat sig att kommissionen på grundval av de första utkasten kommit med mycket viktiga löften .
Vi krävde en föreskrift för " angivare " , och en sådan har kommit .
Parlamentet ville ha en åtskillnad mellan ekonomistyrning och revisionsfunktioner .
Den har vi redan uppnått .
Parlamentet kräver en uppförandekod för kommissionärer och kabinett .
Även det har vi fått .
Parlamentet bad kommissionen att avstå från sina överdrivna förmåner .
Även detta har de gjort .
Samtidigt har kommissionen förpliktigat sig att samarbeta med parlamentet på området SEM-2000 .
Man kommer också att se över kontoren för tekniskt bistånd för att vidta grundläggande förändringar .
Detta är några goda första steg som visar att , om parlamentet så vill , förändringar inte bara är möjliga utan också snabbt kan omsättas i handling .
Vi vill dock ännu mer .
Kommissionen måste nu komma med ett ambitiöst och långtgående reformprogram .
Det är inte bara nödvändigt för en oklanderlig offentlig förvaltning ; det är en conditio sine qua non för att återställa förtroendet hos medborgarna i Europa .
Vi kräver nu tydliga löften av Europeiska kommissionen på följande punkter .
För det första måste parlamentet få fullständig tillgång till kommissionens samtliga handlingar .
Detta står visserligen i motsats till att vi internt snabbt måste nå en uppgörelse för att kunna garantera sekretessen för känsliga dokument .
I samband med inhämtande av information skulle jag vilja göra kommissionen uppmärksam på att vi är mycket oroliga över de preliminära planer som föreligger om allmänhetens tillgång till handlingar .
Om det aktuella utkastet kommer att gå igenom är det ett oerhört steg tillbaka jämfört med i dag .
Det måste bli slut på en situation där finansiellt starka organisationer med representanter i Bryssel kan komma åt information men inte de vanliga medborgarna .
Det får inte heller vara så att en offentlig institution innehar copyright till offentliga handlingar .
Vidare vill vi ha tydliga arbetsbeskrivningar för varje europatjänsteman så att en tjänsteman har dessa samvetsskäl och lättare kan opponera sig mot uppdrag som är oetiska eller olagliga .
Vidare måste det vara så att när revisionsrätten upptäcker att en brist uppträder inte bara ett år utan två år efter varandra bär förvaltningen ansvar för detta , och sådant skall även kunna gå ut över en karriärplanering .
Slutligen måste vi naturligtvis också ha ett bättre samarbete mellan Europeiska revisionsrätten och dess nationella motparter .
Parlamentet kräver också av kommissionen att den den 31 mars i år kommer med en första skiss för reformeringen av den externa biståndspolitiken .
Det får inte längre vara så att Europa visserligen är en ekonomisk makt men att vi inte har något politiskt inflytande därför att vi , när det kommer till kritan , inte kan erbjuda någon effektiv hjälp till områden som verkligen är i behov av sådan .
Som exempel på detta nämner jag Gaza .
Det är oacceptabelt att kommissionen färdigställde ett sjukhus 1996 och att det ända fram till den dag som i dag är inte har legat en enda patient i det .
Herr talman !
Sedan 1996 har ansvarsfriheten fått en tung politisk betydelse .
Det är ett av de starkaste maktmedlen som parlamentet har , och därför måste det användas med försiktighet .
Därför kommer vi med all sannolikhet att bevilja ansvarsfrihet i morgon .
Vi avhänder oss dock inte detta vapen utan att också placera ut en tidsinställd bomb .
Ansvarsfriheten för 1999 kommer nämligen att beviljas först när alla de ekonomiska oegentligheter som revisionsrätten upptäckt har lösts .
Slutligen , denna ansvarsfrihetsrapport riktar sig naturligtvis också till kommissionen .
Men det hindrar inte att också Europaparlamentet måste får ordning på torpet internt .
Så länge vi inte har någon stadga är vi inte trovärdiga som unionens reformeringsmotor .
Reformerna av de europeiska institutionerna är ett nödvändigt villkor för att kunna bygga vidare på Europa .
Det enda sättet att få ett handlingskraftigt och rättvist Europa är att också se till att det är öppet och demokratiskt .
Alla institutioner måste nu slå sig ihop för att tillsammans arbeta för ett sådant Europa . .
( EN ) Herr talman !
Utskottet för industrifrågor bestämde sig för att upprätta ett betänkande om ansvarsfrihet för 1997 trots att vi inte särskilt har ombetts att göra det .
Vi gjorde detta eftersom vi tyckte att vi borde inleda denna mandatperiod på det sätt vi har för avsikt att fortsätta den , det vill säga genom att se till att vi tar väl hand om skattebetalarnas pengar i Europa .
Under vårt arbete på detta betänkande stod det klart att det finns kvarhängande problem inom de utgiftssektorer som ligger i vår budget .
De är inte unika för 1997 och verkar ha två röda trådar .
Den första är kommissionens tendens att ge sig in på mycket ambitiösa program , särskilt i tredje världen , utan att tillräckligt ha utvärderat de praktiska detaljerna kring genomförandet och utan ordentlig resurstilldelning .
Den andra gäller allvarliga administrativa brister hos kommissionen , särskilt vad beträffar samordningen mellan avdelningar och hanteringen av externa kontakter .
Jag vet att alla institutioner har del i ansvaret för kommissionens ökade arbetsbörda och för en del av resursbristen .
Det kan inte ursäkta allt det vi har stött på .
Europas medborgare förväntar sig att de europeiska institutionerna administreras ordentligt och det gör de rätt i .
Det är därför jag vill upprepa min kollegas kommentarer om vikten av den reformprocess som herrar Prodi och Kinnock har lovat Europas folk .
Att döma av det jag har sett av reformprocessen ser det bra ut .
Jag såg några av Kinnocks papper i dag och jag hörde en del av det han hade att säga .
Jag är full av tillförsikt om att vi och Europas politiker kommer att få den slags reform vi behöver om vi stöder honom .
Men vi behöver denna reformprocess .
Många av de generella punkter som tas upp i vårt utskotts betänkande omfattas av van der Laans betänkande .
Det är ett utmärkt betänkande och vi bör alla gratulera henne till det .
Jag tycker att man verkar ha hittat alla de ömma punkterna utan att betänkandet bara blir en uppsättning detaljer , som några av de gamla betänkandena .
De grupperas samman och detta är mycket viktigt .
Jag skulle vilja fästa er uppmärksamhet på två frågor .
Den ena är kärnkraftssäkerhet i Östeuropa .
Vi måste få ordning på detta .
Den oberoende expertkommittén sade att kommissionen inte skötte detta ordentligt .
Vi måste råda bot på detta .
Den andra punkten gäller granskningsmekanismer .
Vi behöver ha material från kommissionen som vi kan använda som hjälp vid granskningen av utgifterna .
Vi behöver ordentlig information som lämnas på rätt sätt och vi måste alla ta hela denna process mycket mer på allvar än vi har gjort hittills .
Den har betraktats som en byråkratisk process som skulle göras så snabbt som möjligt med så liten tidsåtgång som möjligt .
Jag hoppas att kollegerna i denna kammare kommer att stödja skälen för ansvarsfrihet för 1997 och att samtidigt kommissionen kommer att driva på reformprocessen som borde ha genomförts för länge sedan .
Det är enda sättet att skapa en ny kultur i kommissionen och samtidigt återställa allmänhetens förtroende .
Herr talman , kära kolleger !
Parlamentet måste nu fatta beslut om den ansvarsfrihet som den 4 maj förra året förvägrades kommissionen för budgetåret 1997 .
Mot denna för EU verkligt historiska bakgrund måste vi därför fråga oss : Vilka ändringar har skett ?
Vad har förbättrats ?
Vad skulle i dag försvara att man beviljar ansvarsfrihet ?
För det första har vi - i varje fall delvis - en ny kommission .
Vi har fått en mängd avsiktsförklaringar och tillkännagivanden om reformer , alltsammans föga konkretiserat .
Hittills bortser man från skapandet av en uppförandekod för kommissionsledamöter och kabinett .
Jag har också under förmiddagen tagit del av Schreyers utläggningar om överklagandet mot de båda bankerna och stödet för att skapa ett straffrättsligt skydd för EU : s ekonomiska intressen .
Också detta är positiva tecken .
Men man måste medge att de inte kostar kommissionen särskilt mycket .
Kommissionen har varslat om att man skall lägga fram reformprogrammet till februari 2000 .
Nu är tillkännagivanden och avsiktsförklaringar en sak , och genomförandet av givna löften en annan .
Kommissionens ansträngningar kan man emellertid bara bedöma med hjälp av konkreta resultat , eftersom man bara på så vis kan rätta till den enorma brist på förtroende bland medborgarna som EU har drabbats av på grund av inkonsekvenser och manipulationer .
Den summering som vi alltså kan göra sedan i maj 1999 talar inte på något övertygande sätt för ett beslut om ansvarsfrihet .
Om kommissionen trots detta medges ansvarsfrihet för budgeten 1997 så sker det genom att vi garanterar den ytterligare ett stort förskott av förtroende .
Huruvida våra medborgare , med tanke på de svåra överträdelser som begicks av den gamla kommissionen och som naturligtvis betungar den nya kommissionen , över huvud taget kan uppbringa någon förståelse för ett sådant förnyat förtroendeförskott från den demokratiskt valda kontrollinstansen , parlamentet , är en helt annan sak .
Härtill kommer , och det är ändå viktigt för det allmänna intryck som befolkningen får , att revisionsrätten hittills - så vitt jag vet - ännu inte kunnat avge någon positiv revisionsförklaring sedan detta instrument infördes .
Jag förespråkar likväl ansvarsfrihet för 1997 och ber också kollegerna om ett positivt beslut , eftersom man därigenom tar ett tydligt steg och visar att man börjar på nytt , och även ger den nuvarande kommissionen en synlig chans att börja på nytt och få bukt med det erkänt svåra arvet .
Det betyder å andra sidan att alla oriktigheter och bedrägerier även i fortsättningen måste iakttas och klaras upp fullständigt .
Om kommissionen nu medges ansvarsfrihet för år 1997 får detta inte på något sätt uppfattas som om det förgångna är urskuldat eller som ett frikort för framtida bristfällig ekonomisk hushållning .
För när pengar kommer med i spelet tar som bekant vänskapen slut .
Det är ett talesätt som gäller för medborgare såväl som för europeiska institutioner .
Och vänskapen , dvs. i det här fallet förtroendet för tillförlitligheten i de europeiska instansernas arbete , är i dag mer nödvändig än någonsin .
I synnerhet kommer EU : s förestående utvidgning med staterna i Central- och Östeuropa att föra med sig vittgående problem och belastningar även för de inre strukturerna och förvaltningsprocesserna .
En kommission som skakas av ekonomiska skandaler skulle mycket snabbt kunna bli till en lekboll för intressen och mål , som sannerligen inte står på Amsterdamfördragets lista .
Tyvärr har problemen i det förgångna , i synnerhet under det år rapporten gäller , särskilt uppträtt inom de stödområden som i och med utvidgningen tilltar i betydelse , exempelvis strukturfonderna och insatserna från kontoren för tekniskt bistånd .
Detta otillbörliga agerande måste snarast upphöra , eftersom vi inte av de nya stater som ansluter sig kan begära något som vi , de gamla medlemsländerna , inte själva iakttar .
Det är inte heller någon lösning när kommissionen och medlemsstaterna växelvis pekar finger åt varandra och ömsesidigt ger varandra skulden .
Som föredragande för budgeten för 1998 vill jag redan nu meddela att jag under de närmaste veckorna och månaderna kommer att mycket noga iaktta hur och om kommissionen genomför sina reformförslag och hur den utformar sina förbindelser med parlamentet på just detta område .
( Applåder ) Herr talman !
Jag är säker på att kommissionen kommer att bli lättad över att höra att ansvarsfriheten för 1997 troligen inte kommer att få samma konsekvenser som ansvarsfriheten för 1996 vilken , som ni alla är så väl medvetna om , ledde till att Santer-kommissionen tvingades avgå .
Socialistgruppen kommer att rösta för ansvarsfrihet .
Jag är säker på att ni blir lättade av att höra också detta .
Men därmed inte sagt att vi är nöjda , därmed inte sagt att allt är rosenrött .
Det står klart att en radikal omvälvning av kommissionen borde ha gjorts för länge sedan .
Detta betyder emellertid att vi erkänner att de åtgärder man vidtar går i rätt riktning .
Jag vill bara skissera några av de frågor där vi socialister har föreslagit ändringar .
Vi hoppas att dessa kommer att bifallas eftersom de är viktiga på grund av sin inverkan på den kommande reformen .
För det första tjänstemännens immunitet : denna bör upphävas om och när en nationell åklagare så begär .
Vi måste göra det mycket lättare att åtala tjänstemän som har gjort sig skyldiga till bedrägeri och korruption .
Det är avgörande att man noterar att kommissionen allt för ofta har underlåtit att genomföra de reformer som revisionsrätten har rekommenderat .
Det finns skäl till att rättens rapport finns , det finns skäl till vårt svar och det är viktigt att det följs upp .
Jag hörde just att kommissionen kommer att inrätta en arbetsgrupp för revisionsuppföljning .
Så även om vi inte hör någonting mer vet vi att det går åt rätt håll vad beträffar de reformer vi vill ha .
Allt för ofta har vi lagt fram rekommendationer och de har inte lett till någon åtgärd , trots att ni väldigt ofta har sagt att ni skulle handla i enlighet med dem .
Vi vill se denna uppföljning i mycket större utsträckning i framtiden .
Den andra frågan är tillgången till konfidentiella handlingar .
Vi har tidigare haft problem i fråga om vår skyldighet att ta ställning till ansvarsfrihet eftersom vi inte har haft tillgång till de handlingar vi borde ha haft .
Vi inser att även vi har ett ansvar här , att om vi får handlingar måste vi tillse att sekretessbelagda handlingar verkligen förblir sekretessbelagda .
Vi har lagt fram ett ändringsförslag om detta .
En fråga som man hänvisar till i van der Laans betänkande är hela frågan om sjukhuset i Gaza .
Situationen där är helt oacceptabel .
Vi kommer inte att tolerera den mycket längre och vi vill att man omedelbart agerar i denna fråga .
Jag skulle vilja gratulera Lousewies van der Laan .
Vanligtvis bryr jag mig inte om att gratulera människor , men jag tycker att hon har producerat ett mycket övertygande betänkande och förtjänar vårt tack .
Herr talman , kolleger , fru kommissionär !
Låt oss vara ärliga ; vi befinner oss i en något märklig situation .
Vi diskuterar ansvarsfrihet för ett år som ligger bakom oss , men vi diskuterar också kommissionens ansvar .
Jag vill ta upp de problem som fortfarande ligger i skyhöga travar på vårt bord .
Bedömningen i fråga om att bevilja ansvarsfrihet eller inte hänger också i viss mån samman med var man lägger den största tonvikten .
Det handlar om en kommission som inte längre sitter kvar .
Det är en ny kommission .
Då är det logiskt att bevilja ansvarsfrihet , för vad kan den nuvarande kommissionären förebrås för när det handlar om året 1997 ?
De problem som är aktuella finns fortfarande kvar , och då börjar man att tvivla .
Vi måste nu fatta ett beslut om kommissionens goda föresatser , men det föreligger fortfarande ingen strukturerad översikt över dessa goda föresatser .
Kinnock kommer med sitt förslag nästa månad .
Det väntar vi allesammans med spänning på , men vi har ännu inte den kunskapen när vi nu måste fatta beslut om ansvarsfrihet .
Det är tydligen ett dilemma som föredraganden också har brottats med .
Detta dilemma är ännu mer vidsträckt än de områden som jag nämnde .
Det handlar till exempel om kommissionens löften .
De ser i sig bra ut .
Jag har läst ett antal av Kinnocks dokument , och de har vi fullt förtroende för .
Men jag ger två exempel på varför det inte är självklart att de goda föresatser som kommissionen nu gett uttryck för kommer att leda till ett gott resultat .
Offentligheten , sekretessbelagda handlingar .
Detta togs också upp av föregående talare .
Det cirkulerar nu ett dokument , inte på låg nivå utan på hög nivå i kommissionen , varvid offentligheten för dokument inte utökas utan helt enkelt upphävs .
Ett exempel på att ett vackert löfte inte automatiskt kommer att leda till ett gott resultat .
Det gäller också för " angivarna " .
Kinnock har också ägnat dem några vackra ord , men samtidigt är det fullständigt otydligt , just nu när vi skall fatta beslut om detta , vad som till exempel händer med " angivare " som inte får någon chans internt utan som vill gå ut , till pressen , till parlamentet .
Det har fortfarande inte kommit något svar på den sortens avgörande frågor på det området .
Det råder således tvivel , just nu när vi skall fatta beslut om detta , om dessa löften från kommissionen är tillräckligt kraftfulla .
Detta gäller också till exempel för de mycket konkreta projekt som utskottet för industrifrågor har tagit upp .
Jag anser att kommissionen och Kinnock måste komma med goda föresatser , med goda planer för personalpolitiken , för den ekonomiska förvaltningen , men varje kommissionär som nu är ansvarig för ett område med allvarliga brister i det förflutna måste komma med goda planer för att förbättra situationen och inte med allmänna vackra förslag .
För närvarande har vår grupp fortfarande förbarmande , tålamod med kommissionen eftersom den inte kan ställas till ansvar för många felaktigheter ur det förflutna , men detta tålamod är inte obegränsat .
Det måste finnas tydliga framsteg i sikte .
För närvarande förlitar vi oss på att kommissionen kommer med dessa goda förslag , men detta förtroende är inte automatiskt .
Slutligen , herr talman , ansvarsfriheten 1996 var början till slutet för den förra kommissionen .
Jag uttalar förhoppningen , men ännu starkare , jag vill egentligen kräva av den nuvarande kommissionen att ansvarsbefrielsen 1997 är inledningen till en verklig reformering av den ekonomiska politiken från kommissionens sida , för annars kommer denna ansvarsbefrielse inte att ha varit till någon nytta .
När man bedömer frågan om ansvarsfrihet för kommissionen , måste avgörandet grundas på vad som faktiskt hände under det aktuella budgetåret , i detta fall under år 1997 .
I vår grupp har vi svårt att se att den ekonomiska förvaltningen för år 1997 på något avgörande sätt var bättre än den för år 1996 .
Det året röstade vi mot ansvarsfrihet .
I konsekvens med detta kommer vi att rösta mot ansvarsfrihet även för år 1997 .
Vi menar att denna vår bild bekräftas av revisionsrättens granskning .
Det är både bra och nödvändigt att reformer har utlovats .
Ännu så länge återstår det dock att infria de löften som givits , inte minst vad gäller öppenhet .
Vi kommer därför att rösta för de krav på reformer som framförs i resolutionen , men mot att ansvarsfrihet beviljas .
Herr talman !
För det första har jag bara positiva ord att säga om van der Laans mycket väl utförda arbete i samband med detta betänkande .
Gruppen Unionen för nationernas Europa kan inte rösta för ett godkännande av räkenskaperna för budgetåret 1997 .
Betänkandet om s.k. ansvarsfrihet innehåller en omfattande och ytterst kritisk genomgång av räkenskaperna .
Vi stöder dessa kritiska anmärkningar och därför måste jag konstatera att det verkar helt absurt mot denna bakgrund att acceptera ett godkännande .
Det har inte varit möjligt för revisionsrätten att avge en revisionsförklaring om att de dispositioner som räkenskaperna omfattar är lagliga , och vi anser det vara ytterst problematiskt att vi som ledamöter av detta parlament skulle rösta för räkenskaperna utan att säkert veta om dispositionerna är lagliga .
Majoriteten har beviljat ansvarsfrihet under förutsättning att den nya kommissionen genomför en rad reformer som skall se till att det vi erfarit under den förra kommissionens mandatperiod inte upprepas .
Jag måste återigen säga att det handlar om en högst olycklig sammanblandning av den gamla kommissionens ansvar för budgetåret 1997 och den nya kommissionens ansvar för framtiden .
Vi menar inte att den nya kommissionen under några omständigheter skall ha ansvar för den gamla kommissionens politik .
Vi menar att det är felaktigt att tala om kommissionens ansvar som en institution .
Bristerna fram till 1999 skall skyllas på de som då hade ansvaret och vi har ännu inte möjlighet att se om den nya kommissionen kan göra det bättre .
I och med detta märkliga förfarande tar inte parlamentet chansen att placera ansvaret för dispositionerna under budgetåret 1997 där det hör hemma , dvs. hos den tidigare kommissionen .
Det var 1996 års budget som fällde den tidigare kommissionen och 1997 års budget är precis lika betungande .
Det finns inget skäl till att vi mot denna bakgrund skulle bevilja ansvarsfrihet .
Vad gäller beslutet om avslutningen av räkenskaperna vill vi inte delta i omröstningen och slutligen vad gäller resolutionsförslaget vill vi betona de många korrekta godkännandena och rösta för .
Herr talman !
Beslutet om ansvarsfrihet för budgetåret 1997 har skjutits upp , eftersom den kommission som beslutet vid den tidpunkten gällde hade trätt tillbaka och bara var en expeditionskommission .
I dag föreslås det nu i van der Laans betänkande - som hon har lagt ned mycken flit på , och det bör man tacka henne hjärtligt för - att kommissionen medges ansvarsfrihet för budgetåret 1997 .
Man kan fråga sig varför den nuvarande kommissionen får ansvarsfrihet för hur den förra kommissionens skött sin ekonomi - Camre har just berört detta - framför allt som den förvägrades ansvarsfrihet för år 1996 .
Men så ligger det till .
I och med att den nya kommissionen övertog mandatet är den också ansvarig för både goda och dåliga prestationer i det förflutna .
Eftersom kommissionen till sitt system är ett kollegium och endast kan medges ansvarsfrihet i sin helhet , respektive kan få den uppskjuten eller förvägrad , spelar det inte heller längre någon roll att fyra förutvarande kommissionärer hörde till den tidigare kommissionen som hittills inte medgivits ansvarsfrihet , och nu åter är ledamöter i denna institution .
Denna fråga skulle ha behövt ställas när den nya kommissionen tillsattes .
Om parlamentet denna vecka röstar för budgetkontrollutskottets förslag och beviljar ansvarsfrihet , får kommissionen inte förstå detta som en check in blanko .
Ty enligt min åsikt är den tredje delen i van der Laans betänkande den viktigaste , nämligen resolutionsförslaget .
De villkor som samlats under åtta rubriker är väsentliga beståndsdelar av ansvarsfriheten , och vårt beslut utgår från att de uppfylls .
Under processen med beviljande av ansvarsfrihet för åren därefter - 1998 är redan påbörjat - kommer parlamentet att mycket noga få lov att undersöka om det inte alltför snabbt gett kommissionen ett förtroendeförskott för år 1997 .
Det kommer genast att visa sig , när kommissionen lägger fram sitt reformprogram .
Huruvida det då finns någon effektivitet , öppenhet och ansvar , liksom en uttalad informationsvilja gentemot den myndighet som beviljar ansvarsfrihet , kommer vi att granska när ansvarsfrihet för budgetåret 1998 skall beviljas .
Herr talman !
Kollegan van der Laan rekommenderar att man beviljar ansvarsfrihet för budgetåret 1997 , och det uppfattar vi som en vänlig gest gentemot den nya kommissionen , så som föregående talare också har sagt .
Denna ansvarsfrihet medges under förutsättning att kommissionen företar långtgående reformer står det i punkt 1 i resolutionen .
Men den som tror att världen efter avvisandet av ansvarsfrihet för 1996 nu åter är i sin ordning när man medger ansvarsfrihet för år 1997 , har fått saken om bakfoten !
Jag anser att framför allt den frågan är obesvarad , hur långt den nya kommissionen faktiskt är beredd att underkasta sig och sina tjänstemän en kontroll från parlamentets och rättsväsendets sida .
Ett exempel : En av de första frågorna som vi konfronterades med när vi just hade konstituerat oss i budgetkontrollutskottet var det s.k.
Fléchard-fallet , alltså bedrägerier i samband med export av smör till dåvarande Sovjetunionen i början av 90-talet .
Den 7 januari 1994 beslutade höga tjänstemän i kommissionen att efterskänka företaget i fråga det straff det egentligen skulle ha haft , vilket rörde ett belopp om närmare 18 miljoner euro .
Detta innebar att man verkligen överträdde gällande gemenskapsregler .
Vi fick reda på det först genom ett anonymt brev i slutet av 1998 .
Allt jag hittills hört av ledamöter i Prodis kommission kan sammanfattas på så vis att man ändå inte borde fortsätta att gräva i fall som ligger långt tillbaka i tiden , utan hellre se mot framtiden .
Det upprörande här är att generaldirektörer och direktörer , som på sin tid var delaktiga , oskyldigt förklarar för en att protokollet från det avgörande sammanträdet den 7 januari 1994 tyvärr försvunnit på oförklarligt sätt .
Det sägs ha funnits inte bara ett exemplar av det , utan flera .
Varje deltagare skulle ha fått ett exemplar , men alla vore tyvärr omöjliga att återfinna , alla !
När man får höra detta kan man inte längre säga : Låt oss glömma det !
Detta är en händelse som måste finnas med på listan över interna fall som bör undersökas av OLAF , men som såvitt jag vet fortfarande inte finns med där .
Men detta hör också till de händelser som borde meddelas de ansvariga rättsliga myndigheterna , ty när allt kommer omkring är det inte något gentlemannabrott när man ser till att underlag och protokoll försvinner , utan uttryckligen straffbelagt i artikel 241 i den belgiska strafflagstiftningen .
Jag vill bara säga att vi inom ramen för ansvarsfrihetsförfarandet för budgetåret 1998 säkert kommer tillbaka till detta .
Herr talman !
Vi minns alla att parlamentet beslöt att skjuta upp ansvarsfriheten för budgetåret 1997 i avvaktan på åtaganden från den nya Europeiska kommissionen om interna reformer .
Som svar på detta har kommissionen gjort olika åtaganden och har helt klart fattat många beslut om reformer .
I rättvisans namn måste man säga att den nye ordföranden Prodi och hans lag verkligen har förbundit sig att genomföra de mekanismer för ekonomisk kontroll detta parlament har lagt fram .
Reformeringen av Europeiska kommissionen måste dock nu ses mot bakgrund av den debatt som kommer att äga rum inför den kommande regeringskonferensen och reformeringen av olika politiska områden och initiativ inom EU .
Dagens EU-fördrag kommer att ändras för att till exempel säkerställa att utvidgningen kan lyckas .
Jag tvivlar inte på att ytterligare reformer av EU : s institutioner kommer att analyseras i denna debatt .
Men ur de små medlemsstaternas perspektiv är det viktigt att Europeiska kommissionen reformeras på ett sätt som säkerställer att små medlemsstater fortfarande är företrädda i kommissionen .
Herr talman !
Nu får kommissionen sin ansvarsfrihet för budgetåret 1997 , men i realiteten förtjänar de den inte .
År 1997 lyder under den gamla kommissionen och därför menar den nya att den inte kan ta på sig ansvaret .
Det är korrekt att genomförandet av budgeten för år 1997 härrör till den gamla kommissionen , men den nya kommissionen har i gengäld åtagit sig att rensa upp efter de gamla skandalerna och jag måste erkänna att jag inte är särskilt imponerad .
Mentaliteten från förr då man skulle sopa allt under mattan och ställa upp för sina vänner , existerar tyvärr alltjämt .
Det finns vissa som menar att vi är bättre betjänta av att begrava gamla synder och börja på ny kula .
Jag anser att vi inte kan börja på ny kula om vi inte först rensar upp ordentligt .
Jag avser här i synnerhet de gamla skandalerna i ECHO .
Det gör mig mycket irriterad att det är så svårt att få ut handlingar om frågan .
Jag är föredragande för ECHO i budgetkontrollutskottet och det kommer att bli mycket svårt för mig att utföra mitt arbete om inte kommissionen ger mig den nödvändiga informationen .
Utifrån ser det ut som om kommissionen har något att dölja .
Mina undersökningar tyder dessvärre också på att så skulle kunna vara fallet .
Kommissionen lägger inte alla kort på bordet och återupptar alltså sin hävdvunna praxis .
Det var denna praxis som ledde fram till kommissionens fall .
Jag kan därför fullständigt stödja uppmaningen att parlamentet skall ha tillgång till alla handlingar .
I annat fall kan vi inte utföra vårt arbete .
Herr talman , fru föredragande , mina damer och herrar ledamöter !
Jag hoppas att jag kan besvara frågan med ja om vi förtjänar att beviljas ansvarsfrihet .
Tillsammans med revisionsrättens rapport utgör ju ansvarsfrihetsförfarandet när det gäller budgeten den information skattebetalarna erhåller om huruvida och i vilken utsträckning budgetmedel har använts på ett sparsamt sätt och i enlighet med de politiska prioriteringarna , var fel har begåtts , men framför allt också vilka åtgärder som vidtagits med anledning av det .
Att förfarandet med ansvarsfrihet inte betraktas som rutin av Europaparlamentet , utan behandlas mycket noga , det känner allmänheten till , och det vet också kommissionen sedan i fjol , när ansvarsfrihet förvägrades , vilket ledde till att den gamla kommissionen avgick .
Med dagens debatt om ansvarsfrihet för budgetåret 1997 går därför en lång process mot sitt slut .
Den omfattade nästan alla viktiga frågor som kommissionen i vidaste bemärkelse ägnar sig åt .
Van der Laans betänkande berör alla dessa instrument .
Betänkandet är mycket ambitiöst .
Det koncentreras på de reformsteg som inletts , och framför allt på dem som måste påbörjas .
Kommissionen delar föredragandens ambitiösa inställning .
Jag vill gratulera er , fru van der Laan , till detta verkligen mycket ambitiösa betänkande .
Jag vill nu gå in litet närmare på några punkter i betänkandet .
För det första på frågan som med all rätt intar en mycket framskjuten ställning , nämligen frågan om användning av externa resurser för vissa uppgifter .
Vi har diskuterat detta mycket utförligt i utskottet , även inom ramen för budgetförfarandet för år 2000 .
Kommissionen har lovat parlamentet att mycket snart vidta åtgärder här .
Vad gäller kontoren för tekniskt bistånd spelar utrikespolitiken den största rollen .
Min kollega Chris Patten inrättade tillsammans med de andra kommissionärerna , som är ansvariga för utrikespolitiken , redan i slutet av förra året en Review-grupp , som mycket snart skall gå igenom nuvarande kontor för tekniskt bistånd med tanke på deras uppgifter , och granska vilka som i framtiden bör få en annan form .
Gruppen har föresatt sig att kort efter att hela reformpaketet lagts fram också komma med speciella förslag för detta utrikespolitiska område .
Det kommer troligen inte att bli möjligt för kommissionen att redan den 31 mars lägga fram ett detaljerat förslag om denna speciella punkt , men , hoppas vi , mycket snart därefter .
Ni hade hänvisat till totalkonceptet i ert betänkande .
Detta totalkoncept är en beståndsdel i reformpaketet .
Men jag ville också nämna att konkreta åtgärder förbereds för detta utrikespolitiska område - även i enlighet med Bourlanges betänkande .
Andra krav i betänkandet syftar till att öka insynen .
Även här vill jag försäkra att ni där berör en av de reformer som kommissionen syftar till .
Den vill vara en öppen kommission , som möjligen inskränker informationen gentemot er kammare när det gäller intressen som måste skyddas .
Jag hyser tillförsikt för att dessa frågor kommer att kunna regleras i det interinstitutionella avtalet .
Kommissionen kommer även att förbättra informationsnivån på sina räkenskaper , utöver existerande rättsliga förpliktelser , som krävs av er och revisionsrätten .
Redan vid debatten om revisionsrättens rapport lovade jag att jag tar upp denna punkt , som också finns med här i betänkandet , nämligen att göra en systematisk follow-up , eftersom jag anser att det är nödvändigt .
Kommissionen har på mitt förslag redan beslutat ge revisorerna i uppdrag att redan i bokföringen för år 1999 ta hänsyn till revisionsrättens kritik , nämligen att i bokföringen föra förskottsbetalningar separat , så att denna information finns till hands .
Bekämpningen av bedrägerier skall förstärkas ytterligare .
Vi har också redan under förmiddagen kort diskuterat OLAF .
Den i budgeten 2000 upptagna ökningen av personalen vill jag nämna än en gång .
Fru Stauner , det överklagande jag nämnde i förmiddags har ju inte bara utlovats , utan redan lämnats in .
Jag tror att detta också visar att kommissionen inte är beredd att acceptera att vissa institutioner vill undandra sig dessa bestämmelser som beslutats av parlamentet och rådet , utan de sträcker sig ju till alla institutioner inom Europeiska gemenskapen .
Slutligen kräver ni också en förbättrad dialog , mer dialog med medlemsstaterna om nödvändiga förbättringar när man beslutar om gemenskapsmedel .
Även här stöder jag era krav och kommer att hålla ögonen på att det genomförs i de fall där kommissionen berörs .
Beträffande frågorna om sjukhuset i Gaza och det palestinska parlamentet kan jag meddela er att sjukhuset i Gaza kommer att vara öppet och stå till förfogande för läkarbesök från och med den 15 juli , och för sjukhusvistelser från och med den 15 oktober 2000 .
För det andra kommer kommissionen att till den 31 mars informera Europaparlamentet om de framsteg som görs vad gäller sjukhuset och val av de consultants , som skall förbereda handlingarna för anbudsförfarandet för byggandet av det palestinska parlamentet .
Alla reformåtgärder som jag har berört är delar av ett totalkoncept .
Min kollega Kinnock kommer att lägga fram kommissionens helhetskoncept för er , och tala om de politiska prioriteringarna under denna mandatperiod , liksom om detaljkonceptet , med avseende på en konkret och framför allt kontrollerbar och förståelig tidsplanering .
Genomförandet av dessa planer skall i sin helhet göra Europeiska unionen och dess institutioner mer slagkraftiga och öppna .
Det är parlamentets uppgift , i synnerhet inom ramen för förfarandet beträffande ansvarsfrihet , att kontrollera kommissionens verksamhet .
Kommissionen är sannerligen medveten om hur konkret och exakt Europaparlamentet genomför denna kontroll .
Jag är desto gladare över att de inledda reformåtgärderna bedöms positivt av er , och att ni är beredda att besluta om ansvarsfrihet för budgetåret 1997 .
Tack så mycket , kommissionär Schreyer !
Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
 
Åtgärder att vidta med anledning av den oberoende expertkommitténs andra rapport Nästa punkt på föredragningslistan är betänkande ( A5-0001 / 2000 ) av van Hulten för budgetkontrollutskottet om åtgärder att vidta med anledning av den oberoende expertkommitténs andra rapport om reformering av kommissionen . .
( EN ) Herr talman !
Vid den här tiden förra året inrättade Europaparlamentet en oberoende expertkommitté med Middelhoek som ordförande , som skulle granska anklagelser om bedrägeri , nepotism och korruption i Europeiska kommissionen .
15 mars offentliggjorde kommittén sin första rapport med slutsatsen att : " Det börjar bli svårt att hitta någon som har någon som helst ansvarskänsla " .
Bara några timmar efter det att rapporten hade framlagts tillkännagav ordförande Santer att hela hans kollegium avgick .
Avgången markerade slutet på en bitter kamp mellan ett allt mer självsäkert parlament och en kommission som var befläckad av skandalanklagelserna .
Sedan dess har situationen i Bryssel förändrats till oigenkännelighet .
Ett nytt parlament med en ny vigör har valts och en ny kommission tillsatts .
När den nominerade ordföranden Prodi talade i denna kammare 21 juli förband han sig att beakta den andra rapporten från den oberoende expertkommittén för reformering av kommissionen fullt ut .
Denna innehåller 90 detaljerade rekommendationer och det är den vi diskuterar i dag .
Den nya kommissionen har redan tagit viktiga steg bort från sitt gamla sätt att fungera .
En uppförandekod för kommissionärer och deras kabinett har antagits .
Som en symbolisk men betydelsefull gest har kommissionärerna frivilligt avstått från sin rätt till skattefria inköp av alkohol , tobak , bensin och konsumentvaror .
Nya regler har tagits fram och förverkligats vad beträffar hur högre tjänstemän utses .
Antalet avdelningar har minskats .
Enligt min mening har kommissionen visat ett tydligt engagemang utan tidigare motstycke för förändring och detta skall de ha en eloge för .
Det övergripande syftet med reformerna måste vara att skapa en stark , ärlig europeisk offentlig sektor som är rustad för att genomföra sina uppgifter på ett effektivt och kompetent sätt , en offentlig sektor där tjänstemännen har medel att genomföra sina uppgifter och hålls fullt ansvariga på alla nivåer , en offentlig sektor som känner igen och belönar det förtjänstfulla och uppmuntrar tjänstemännen att utveckla hela sin potential .
För att uppnå detta måste vi agera på fyra områden .
För det första måste den ekonomiska hanteringen och kontrollen inom kommissionen förbättras .
Ett av de största problemen är att det saknas ett fungerande system för ekonomisk kontroll .
Kommissionens generaldirektorat måste få ett totalansvar för sina egna kostnader , inklusive den ekonomiska kontrollen .
Ett nytt oberoende revisionssystem måste införas .
Generaldirektoraten måste offentliggöra sina egna årsberättelser så att problemområden tydligt kan identifieras och uppställa årliga mål för att minska bedrägerier och regelbrott .
I utbyte för denna större självständighet måste cheferna göras fullt och personligen ansvariga för sitt agerande .
Det är klart att övergången till ett sådant nytt system kommer att ta tid .
Det kommer att krävas förändringar i budgetförordningen och parlamentet måste uttala sig om dessa förändringar .
Men även om kommissionen måste se till att den följer fördraget och budgetförordningen under en övergångsperiod får inte detta bli en ursäkt för att inte göra någonting .
Det finns ett trängande behov av förändringar i dag .
För det andra måste kampen mot bedrägeri , misskötsel och nepotism intensifieras , främst genom att man skapar en kultur där de inte kan frodas .
Detta kräver att kommissionärerna och de högre tjänstemännen statuerar klara exempel och erbjuder lämplig utbildning , och dessutom att de befintliga mekanismerna för att hantera bedrägerier förstärks .
OLAF , kommissionens byrå som skapades tidigare i år , måste sättas under en oberoende europeisk allmän åklagares ledning , vars uppgift skall vara att förbereda åtal i nationella brottmålsdomstolar av kriminella handlingar som begåtts mot unionens ekonomiska intressen av ledamöter och tjänstemän i de europeiska institutionerna .
Ett förslag kan läggas , ett förslag bör läggas , på grundval av artikel 280 i fördraget senast vid halvårsskiftet .
För det tredje måste det europeiska offentliga livet uppfylla högt satta normer .
Den politiska kris som ledde till att kommissionen föll tidigare i år visade tydligt på behovet av otvetydiga uppföranderegler vars efterlevnad kan framtvingas .
Ett antal koder har sedan införts .
De måste utvärderas av parlamentet och bör göras juridiskt bindande .
De europeiska institutionerna bör följa det exempel som ett antal länder har satt , i synnerhet Storbritannien , och tillsätta en kommitté för normer i det offentliga livet med mandat att ge råd om yrkesetik och uppföranderegler inom de europeiska institutionerna .
Uppgiftslämnare som är i god tro måste skyddas .
I slutet av förra året tillkännagav Kinnock nya åtgärder för att skydda uppgiftslämnare .
Dessa måste genomföras utan dröjsmål .
Även om sådana åtgärder aldrig kan bli ett alternativ till en god ledning måste det finnas en säkerhetsventil när någonting går fel .
Det är avgörande att reformerna inte begränsas till kommissionen .
Även parlamentet måste överväga behovet att förbättra sina interna regler , administrativa rutiner och ledningsutövning .
Slutligen måste kommissionens personalpolitik moderniseras .
Den är helt klart inte anpassad till kraven från en modern , multinationell organisation .
Den sociala dialogen har ofta fungerat som en broms för reformer och borde ha setts över för länge sedan .
Det måste bli mer attraktivt att arbeta inom de europeiska institutionerna .
Allt för många unga , nya tjänstemän lämnar sina jobb efter bara några år .
Förtjänster måste erkännas och belönas , specialutbildning måste bli ett sine qua non för befordran till högre befattningar .
Befordringssystemet måste göras rättvisare och ges ökad insyn .
Sist men inte minst måste löne- och förmånspaketet ses över .
Det måste bli flexiblare och visa större ansvar för arbetsmarknadens villkor .
Det måste befrias från vissa av sina mest förlegade beståndsdelar och man måste ta itu med den berättigade kritiken från allmänheten , som inte kan inse varför EU : s tjänstemän skall få utflyttningsbidrag i all oändlighet i ett Europa med öppna gränser eller betala skatter vars nivå ofta ligger långt under nivån i medlemsstaterna .
Kommissionär Kinnock kommer att framlägga sitt meddelande om reformerna i morgon .
Detta meddelande måste innehålla en klar tidtabell .
Med en ny kommission och ett nytt parlament i full gång är incitamentet för reformer starkare än det någonsin har varit och förmodligen någonsin kommer att bli .
Utvidgningen av unionen ligger bara några år framåt i tiden .
Nu är det dags för Europa att göra rent hus och inpränta en ansvarskänsla - som de oberoende experterna kunde ha sagt - hos sina institutioner .
I juni förra året gav väljarna i Europa en tydlig signal om att de är trötta på ändlösa historier om misskötsel och nepotism .
Det finns ett mycket enkelt sätt att handskas med dessa historier .
Låt oss avskaffa misskötsel och nepotism .
Herr talman !
Jag hoppas verkligen att ingen missförstår mig och därför vill jag först av allt säga att jag naturligtvis är för en kamp mot bedrägeriet och att jag med kraft stöder alla lämpliga och nödvändiga reformer .
Detta är en fråga som inte är enkel och som skulle behöva fördjupas betydligt mer , men jag kommer att nöja mig med att bara peka på enstaka punkter , bl.a. för att ni , om möjligt , skall bli medvetna om vad vi talar om .
Experterna kan ge information och upplysningar , formulera uppfattningar och ge råd , men de har inte något politiskt ansvar gentemot sina väljare .
I stället är det politikerna som måste undersöka vad de kan utnyttja i en expertrapport och vad man inte kan tillämpa i sin helhet i en anda av , som det ibland har verkat , självplågeri .
Jag tror - låt mig bara nämna ett par punkter - att när det gäller ledamöterna i detta parlament så är det enbart parlamentet självt som kan agera och ingen annan , för om det inte var så , så skulle Europaparlamentets auktoritet och representativitet allvarligt hotas under de kommande åren och vår institution skulle inte utvecklas så som den borde .
Det är minst lika viktigt att ingen skall kunna vägra lämna ut handlingar till Europaparlamentet och dess utskott .
Moral , disciplin och sekretess när det gäller de frågor som delegeras skall vara något som avgörs av ledamöterna i detta parlament , och inte något som bestäms utifrån av någon annan .
Låt mig understryka att det inte existerar någon europeisk lag , utan ett diversifierat rättssystem i de olika medlemsstaterna .
Vi löper risken att delegera frågor som rör samma brott och som sedan kommer att bestraffas olika .
Jag håller med om att man bör inrätta ett undersökningssystem , men jag är lika djupt övertygad om att man måste ge rätten att försvara sig samma möjligheter och samma ställning .
Jag håller inte med om att man hur enkelt som helst skall kunna göra Europeiska gemenskapens tjänstemän till brottslingar : angiveri är en metod som inte hör hemma i det tredje millenniet .
Avslutningsvis vill jag säga , herr talman , att från detta parlament bör utgå en tydlig signal om demokratiska principer : vi skall genomföra reformer som gör att parlamentet växer och som utvidgar dess befogenheter , inte som gör att det går tillbaka i utvecklingen .
Denna debatt om van Hulthens betänkande avslutar en av de mest traumatiska perioderna för de europeiska institutionerna sedan de skapades 1957 .
Europaparlamentets vägran att bevilja ansvarsfrihet och den definitiva vägran att bevilja ansvarsfrihet för 1996 års budget , den misstroendeförklaring som bordlades i denna kammare av olika skäl för ett år sedan och den första rapporten från den oberoende expertkommittén om reformering av kommissionen som ledde till kommissionärernas massavgång är nu europeiska folksägner .
De av oss som var inblandade i dessa historiska händelser är väl medvetna om att inga av dessa omvälvningar skulle ha skett om vi inte hade agerat med parlamentarisk makt för att kräva förändringar i kommissionens sätt att fungera .
Minns att ministerrådet , som är frånvarande igen denna debattkväll , beviljade ansvarsfrihet för 1997 - inte 1996 - samma dag som kommissionen avgick , 15 mars .
Nu har vi kommit till den andra rapporten från den oberoende expertkommittén , vilken vi redan har haft tillfälle att välkomna och kort debattera i september .
Det viktigaste för oss i PPE är att tillse att allmänhetens förtroende för Europeiska kommissionen återställs .
Ytterligare steg för att bygga ett starkt Europa kommer inte att tjäna någonting till om de europeiska folken uppfattar att det inte finns något lämpligt system för demokratisk kontroll av övernitiska tjänstemän .
Inte under några omständigheter kommer vi att släppa i från oss de landvinningar vi har gjort under de senaste månaderna , vilka vi tror är till gagn för öppenheten och insynen .
Det bekymrar oss därför att se skurarna av tillkännagivanden från kommissionen under de senaste veckorna där kommissionär Kinnock lägger olika policyförslag som skall ingå i en vitbok som snart kommer .
Detta avslöjar en önskan att gå snabbt fram , men det ger också intrycket att kommissionen befinner sig i sändningsläge snarare än i lyssningsläge .
Vår oro förstärks om det rykte som rapporterades för några dagar sedan stämmer - nämligen att kommissionen kraftigt vill begränsa parlamentets tillgång till information .
Detta var när allt kommer omkring en av orsakerna till att den förra kommissionen föll .
Har man inte lärt sig läxan ?
Vetskapen om att ramen för förhållandet mellan Europaparlamentet och Europeiska kommissionen ännu inte är framförhandlad ledde till att vi var oense med föredraganden när vi diskuterade hans betänkande i utskottet .
Vi kunde absolut inte instämma i hans åsikt att det skulle vara förnedrande för parlamentet att ta fram detaljerade instruktioner om vad vi vill att kommissionen skall ta upp i sitt reformpaket .
Ju mindre exakta vi är i våra resolutioner , van Hulthen , ju mer utrymme får kommissionen och era tidigare kolleger i rådet att göra vad de vill .
Vi anser att det stora antalet rekommendationer i den oberoende expertgruppens rapport bör genomföras .
Vi har , för PPE-DE-gruppens räkning , framlagt alla rekommendationerna i expertgruppens rapport för utskottet , och många av dem har nu tagits med i betänkandet vilket helt förändrar van Hulthens betänkande i utskottet .
Vi har framlagt några ändringsförslag som föll i utskottet , särskilt vår önskan att uppförandereglerna skall ses över .
Främst vill vi lägga in hänvisningen till förtjänster och ledarförmåga som ni , herr kommissionär , när vi hade vår utfrågning i september , accepterade skulle innefattas i dessa uppförandekoder , särskilt beträffande tillsättningar och befordran .
När vi ser framåt vet vi att vi befinner oss i början av en lång process av kontinuerlig reformering av Europeiska kommissionen .
Vi vill särskilt se att bilden av kommissionens tjänstemän som hårt arbetande och mycket kompetenta bekräftas av yttervärlden - ett rykte som har fördunklats av ett fåtal individers olämpliga uppträdande .
Herr kommissionär , ni är säkert medveten om varför krisen uppstod eftersom ni var med i den förra kommissionen .
I ett nötskal : programverksamhet bedrevs utan att det fanns tillräckliga personalresurser tillgängliga .
Vi uppmanar er att ta tillfället i akt att fastställa det verkliga bemanningsbehovet för kommissionen på basis av den viktiga verksamhet den ansvarar för .
Vår inställning i budgeten för 2000 var mycket klar i denna fråga .
Vi kommer att vara vaksamma de närmaste fem åren för att säkerställa att de reformer som nu föreslås genomförs fullt ut och vi kommer att stödja ansträngningar att modernisera institutionerna .
Men å andra sidan kommer vi inte att tveka att dra in vårt stöd vad gäller det finansiella eller annat om åtgärder skulle vidtas som inte överensstämmer med den öppenhet kommissionens ordförande Romano Prodi lovade innan han utsågs .
Låt oss hoppas att vi kan undvika institutionella omvälvningar genom att föra en ständig dialog som från början utgår ifrån att parlamentet skall vara en jämställd partner i besluten om reformeringen av kommissionen .
Herr talman !
Jag måste börja med att be om ursäkt för att jag inte kan vara tillnärmelsevis så dramatisk som Elles i min föredragning .
Låt mig först tacka van Hulthen för hans betänkande .
Det är ett utmärkt betänkande .
Det skulle ha varit fel av parlamentet att okritiskt stoppa in varenda rekommendation från ett utomstående organ , för parlamentet bör ha en egen uppfattning om dessa frågor .
Det är rätt att vi har ett fokuserat betänkande , vilket är vad van Hulthen har producerat .
Tillåt mig att uppmana Elles att inte spänna vagnen framför hästen .
Ja , socialisterna förlorade en hel del saker men de har inte gått igenom i plenum än och låt mig varna honom för att de kanske inte gör det i morgon .
Jag skulle vilja tacka kommissionär Kinnock för alla hans ansträngningar hittills .
Han har varit tydlig om att han har förpliktigat sig att genomföra en radikal förändring .
Försöket att skapa och införa ansvar är centralt i detta .
Det är klart att detta måste utvecklas på alla nivåer och att man måste uppfatta behoven på alla nivåer inom kommissionen .
Det står klart att vi behöver en förändring av budgetförordningen .
Detta är viktigt .
Vi måste sätta stopp för att människor skyller ifrån sig på varandra .
När fel uppstår inom kommissionen måste vi ställa någon till ansvar .
Vi måste få försäkringar om att konsekvent underlåtenhet att sköta sina uppgifter skall leda till avsked .
Detta är naturligt på andra håll , men tycks vara ett extremt radikalt förslag när det ställs till kommissionen .
Vi kan inte fortsätta med en situation där inkompetens , misskötsel och bedrägeri kostar de europeiska skattebetalarna pengar och ger dem dålig service .
Jag skall ge er ett exempel på detta .
I revisionsrättens rapport för 1998 kostade en felberäkning av växelkurserna beträffande italienskt vin Europas skattebetalare mellan 8 och 10 miljoner brittiska pund .
Det står klart att detta inte är acceptabelt .
Vad hände med den person som var ansvarig för felräkningen ?
Vi behöver ett system som ger incitament och befordran och denna befordran skall ske på grundval av meriter .
Vi inser att de flesta av tjänstemännen inom kommissionen arbetar extremt hårt .
Men vi inser också att vissa rutiner är föråldrade .
Vi ser fram emot att få läsa kommissionens hela förslag till reform och vi ser fram emot att utarbeta detaljerna jämsides med kommissionen för , trots det Elles just sade , har kommissionären gjort ett åtagande att diskutera det med parlamentet före den 1 mars .
Vi måste också inse att man inte skall kasta sten i glashus .
Europaparlamentet har inte precis varit snövitt i sitt uppträdande under historiens gång .
Vi har långt kvar innan vi är perfekta själva .
Vår egen personalpolitik är förlegad .
Vissa av våra arbetsrutiner behöver reformeras radikalt .
Jag hoppas att Europaparlamentet kommer att hålla fast vid kommissionens rockskört i denna reformprocess .
Vi godkänner förslagen om verksamhetsbudgetering .
Vi inser att detta innebär disciplin från kommissionens tjänstemäns sida och vi inser också att vi har ett ansvar i parlamentet för disciplin när vi talar om negativa prioriteringar .
Låt mig slutligen säga att kommissionen behöver arbeta på sina relationer med allmänheten .
Europas skattebetalare behöver lugnas .
Kommissionens öde , hela Europeiska unionens öde , beror på om denna reform kan genomföras .
Detta är huvudfrågan , att dessa förslag genomförs .
Herr talman !
Jag skulle vilja börja med att framföra mina komplimanger till föredraganden , herr van Hulten , för hans första betänkande .
Jag beundrar honom särskilt för att modet inte svek honom när han drunknade i så många ändringsförslag .
Jag tror att den oberoende expertkommitténs rapport har varit en nyttig rapport , och jag tror också att det är nyttigt för parlamentet - vilket också Morgan sade - att vi också för en gångs skull ber expertis utifrån att se över hur vår administration sköts .
Vi har lagt fram ett ändringsförslag om detta .
Jag skulle vilja understryka ett par av de många punkterna i van Hultens betänkande , det beror inte på hur pass viktiga de är utan det är helt enkelt godtyckligt .
Först och främst anser jag att kommissionen måste ägna mycket större uppmärksamhet åt att bevara dokument på ett betryggande sätt .
Kommissionens arkiv lämnar åtskilligt övrigt att önska .
Vi lade märke till detta när vi skulle undersöka Fléchard-affären som för övrigt inte på långa vägar är utredd ännu .
Konstigt nog hade mycket viktiga dokument försvunnit från kanslierna , till och med från ordförandens , från olika generaldirektorat , och det är helt klart något som inte får förekomma .
Om parlamentet vill göra en ordentlig kontroll måste dessa dokument vara tillgängliga , och jag skulle gärna vilja veta vad kommissionen tänker göra för att förbättra detta .
Sedan något om kontrollen i efterhand , revisionsförklaringen .
Det har också delvis framkommit i van Hultenbetänkandet .
Jag tror att det skulle vara bra om vi började ge rapportsiffror per kategori och per sektor om hur budgeten verkställs .
Nu är det allmänna intrycket att allt i Europa som har med budgeten att göra är dåligt .
Det står klart att vi under de senaste åren sett en förbättringstendens i fråga om jordbruk och en försämrande sådan i fråga om utgifterna för strukturella åtgärder .
Är det acceptabelt ?
Jag skulle vilja föreslå kommissionen att fastställa en deadline för genomförandet av strukturutgifterna .
När vi antar nya medlemsstater får det inte vara så att vi ännu inte bringat ordning i eget hus .
Herr talman , kolleger !
Först och främst vill jag rikta ett tack till kollega van Hulten .
Det är hans första betänkande här i plenum .
Det är värt att gratulera , även om jag naturligtvis beklagar att han inte förklarat detta betänkande på sitt eget modersmål .
Bästa kolleger !
Det är ett betänkande som varit svårt att få till stånd , och kanske kommer det för sent .
Det har enligt min uppfattning framför allt att göra med bråket mellan de två stora grupperna i vårt budgetkontrollutskott .
Låt oss vara ärliga .
Den andra rapporten från den oberoende expertkommittén kom i september .
Nu har det gått ytterligare fyra månader .
Under tiden har van Hulten drunknat i ändringsförslag , mer än 100 ändringsförslag under den första omgången .
Han satte i gång på nytt , skrev om sitt betänkande , tog hänsyn till en stor mängd förslag , men möttes av ytterligare nästan 100 ändringsförslag under den andra omgången .
Allt detta har således lett till , och det är jag litet orolig för , att betänkandet blivit för detaljerat , för omfångsrikt och framlagt för sent .
Dessutom godkände , efter vad jag fått höra , kommissionen alldeles nyligen i dag ett förslag om reformeringen av kommissionen som kommer att skickas runt till olika institutioner för vidare konsultationer och även till vårt parlament hoppas jag .
Skulle Kinnock kanske vilja lyfta på förlåten redan i kväll ?
Kollega van Hulten !
Min grupp av gröna och regionalister kommer inom kort att stödja förslagen under plenum i morgon eftermiddag om att ytterligare förbättra detta betänkande något .
Det ju ingen mening med att ord för ord ta upp de många goda rekommendationerna från den oberoende expertkommittén i ert betänkande .
När vi i morgon således kommer att rösta emot vissa ändringsförslag eller emot vissa punkter är det absolut inte på grund av innehållet , utan i avsikt att göra en mer läsbar helhet av ert betänkande .
I vilket fall som helst måste det stå klart att min grupp naturligtvis fullständigt stöder rekommendationerna från den oberoende expertkommittén .
Hur som helst ser jag fram emot det dokument som godkänts av kommissionen i dag .
Hur som helst ser jag fram emot den vitbok som skall komma inom kort i februari .
Hur som helst måste jag meddela er , herr kommissionär , att både expertkommitténs rapport och van Hultens betänkande kommer att bli riktpunkter för vår grupp , riktpunkter som kommer att tydliggöra för oss om vi , ja eller nej , skall kunna hysa misstroende eller förtroende för kommissionen Prodi .
Som avslutning vill jag bara säga detta .
Precis som i fråga om vitboken om livsmedelssäkerhet som godkändes förra veckan och släpptes till allmänheten och som innehöll en konkret tidsgräns vill vi att detta också skall gälla för den nya vitboken om reformeringen av kommissionen .
Jag tror att detta är nödvändigt eftersom allmänheten ser fram emot förändring , och i vilket fall som helst vill min grupp att en tydlig förändring har förverkligats fram emot slutet av år 2002 .
Herr talman !
Det är bra att detta betänkande har kommit till , men det behövs egentligen mer .
Bedrägeri , dålig förvaltning och svågerpolitik uppstår inte av en slump .
De får den största chansen om den demokratiska kontrollen av penningflödena är ringa .
Via strukturfonderna pumpas en stor del av den europeiska budgeten runt .
Det är meningsfullt endast så länge det handlar om solidaritet där rika medlemsstater bidrar till fattigare medlemsstaters inkomster och utveckling .
Men det förekommer också pengar som pumpas runt och som via Bryssel åter går till samma rika medlemsstater .
Kommuner och regionala myndigheter ser detta som sina egna pengar , men det enda sättet för dem att få dessa pengar är genom att lägga mycket pengar och arbetsinsatser på lobbyverksamhet och förhandlingar .
Efter varje oavsiktlig användning av dessa pengar , och självfallet efter bedrägeri , ljuder ropet på ännu strängare kontroll .
Inte ens den allra strängaste kontroll kan lösa detta problem .
Den kommer på sin höjd att leda till mer byråkrati och mindre utrymme för den lokala demokratin att vinna inflytande och mindre utrymme för medinflytande för befolkningen över val av projekt och deras innehåll .
Det är bättre om dessa pengar slussas direkt från de nationella myndigheterna till de lägre myndigheterna utan att ta omvägen över Europa .
Vi måste någon gång under de kommande åren tänka över möjligheten att ersätta strukturfonderna med en utjämningsfond som är begränsad till budgetstöd för medlemsstater eller deras delstater med en låg inkomst per capita hos befolkningen .
Det är förmodligen den enda vägen för att nå fram till mindre bedrägeri , mindre overhead-kostnader , mer öppenhet och mer demokrati .
Herr talman !
Det har fortfarande inte gått ett år och det är redan en uppenbar skillnad mellan det sätt på vilket parlamentet behandlar det första och det andra betänkandet .
Det första betänkandet gavs omfattande publicitet , det diskuterades högtidligt och utnyttjades därefter , tillsammans med den polemik och de läckor till pressen som föregick det , till att massakrera kommissionens ordförande och därefter de flesta av kommissionärerna , trots att de inte hade något att göra med bedrägerier , tjänstefel och nepotism .
När man nu läser det som hände för knappt ett år sedan verkar det tydligt att det betänkandet skulle kunna användas till vad som helst utom att skapa klarhet eller genomföra reformer , som man hävdar i dag .
På samma sätt är det sant att detta andra betänkande , som i stället skulle kunna lägga fram betydligt konkretare uppgifter , beställdes i det uttalade syftet att inte behandla specifika fall , varför det knappast är intressant att följa upp de olagligheter som nämns .
Det intresserar inte de stora grupperna i detta parlament , och inte heller de flesta av de fackföreningar som i ord anstränger sig att försvara den europeiska förvaltningen , men som i själva verket bara är intresserade av att skydda sina egna medlemmar , och att därvid på ett diskutabelt vis använder de omfattande maktbefogenheter de tilldelats .
Fackföreningsrepresentanter finns det i disciplinråden och i kommittén för tjänsteföreskrifterna , vilket gör det omöjligt att avlägsna de felande tjänstemännen eller att ändra på tjänsteföreskrifterna .
Fackföreningsrepresentanter sitter också , obegripligt nog , i urvalskommittéerna , och jag skulle inte bli förvånad om inte företrädare för fackföreningarna också ingår i OLAF , vilket gravt skulle skada denna institution som åtminstone formellt borde kunna ge garantier om att stå fri från de olika parterna .
Jag förstår med andra ord varför vi träffas vid denna tidpunkt , som i regel är avsedd för annat och inte för debatt , diskussion och information .
Herr talman !
I van Hultenbetänkandet understryker parlamentet den bittra nödvändigheten av en grundlig reformering av den ekonomiska förvaltningen .
Kontrollen av utgifterna måste förbättras kraftigt , såväl hos kommissionen som i medlemsstaterna .
I detta syfte måste även Europeiska revisionsrätten och de nationella revisionsrätterna samarbeta bättre .
Vidare finns det behov av föreskrifter för uppgiftslämnare .
Alla dessa rekommendationer stöder vi helhjärtat .
Men jag har några randanmärkningar .
En av den oberoende expertkommitténs slutsatser är att den nuvarande rättsliga ramen för bekämpning av bedrägeri är osammanhängande och ofullständig , vilket är till nackdel för Europeiska unionen .
I vilken riktning skall vi ta itu med detta ?
Inte genom att frånta medlemsstaterna rättsliga befogenheter och överföra dem till en europeisk åklagarmyndighet .
Någonting sådant förutsätter en europeisk straffrätt , och den finns över huvud taget inte .
Detta berör dessutom kärnan i medlemsstaternas suveränitet .
Därför måste vi söka efter lösningen i ett bättre samarbete mellan medlemsstaterna på det rättsliga området .
Samordningen av detta skulle kunna ske genom en sorts europeisk allmän åklagare .
Denne får inte själv inleda åtal , utan överlämnar brottsärenden till de nationella rättsliga myndigheterna .
Rapporten från den oberoende expertkommittén har också haft ett sanningens ord att säga rådet och parlamentet .
Rådet måste till exempel tillerkänna förfarandet för ansvarsfrihet för kommissionen betydligt större vikt .
I lika hög grad måste parlamentet ta upp den kastade handsken .
Det är verkligen på tiden att det nu kommer en stadga för ledamöter och en resekostnadsersättning på grundval av de verkliga utgifterna .
Detta väcker frågan om parlamentet verkligen är berett att ta sig ur dödläget .
Denna vecka har Rothleys yttrande diskuterats i utskottet för rättsliga frågor , och ingenting i detta visar på någon sådan beredvillighet .
Herr talman !
När det gäller er egen reform , är kommissionen i knipa .
Efter de händelser som ledde till att den tidigare kommissionen avgick , finns det en enorm förväntan .
Jag får ibland intrycket att förslagen även här i kammaren får större bifall , ju mer radikala de låter .
Å andra sidan kan man inte enbart med ett par penndrag ändra på förhållandena från i dag till i morgon , och svårigheterna börjar så snart det gäller genomförandet , så snart man skall tala om detaljer .
Det är möjligen förklaringen till varför vi också i budgetkontrollutskottet haft fler svårigheter än väntat .
Trots detta kan resultatet som det nu föreligger ses som beaktansvärt , och jag vill uttryckligen tacka kollegan van Hulten för hans arbete med detta betänkande .
Om detta betänkande nu inte än en gång urvattnas genom att man antar ändringsförslag , ger vi därmed kommissionen på några avgörande punkter klara och otvetydiga uppgifter .
Låt mig börja med den viktigaste uppgiften .
Vi vill inte avskaffa ekonomistyrningen .
Det måste även i fortsättningen vara möjligt för styrekonomen att göra en granskning innan ekonomiska åtaganden eller betalningar genomförs , inte i alla enskilda fall , men alltid där det finns osäkerhet eller risker .
Här ger kommissionen fel signaler , till exempel när man döper om Generaldirektoratet för ekonomistyrning till Generaldirektorat för revision .
Kommissionens organisationsschema går väl lätt att ändra , men det blir svårare när kommissionen angriper lagtexterna , i synnerhet budgetförordningen .
Jag har inte räknat efter så noga , men gemenskapens budgetförordning och de dithörande genomförandebestämmelserna talar på nästan 100 olika ställen om styrekonomen , hans oberoende och de uppgifter han har .
Detta kan inte ignoreras eller kringgås , inte heller med s.k. soft law , som det en gång antyddes under ett sammanträde med vårt utskott .
Oberoende av sådana rättsliga överväganden vore det också med tanke på sakens natur ett oförlåtligt fel att avskaffa ekonomistyrningen i dess klassiska bemärkelse just i det ögonblick , när de i kommissionen som är ansvariga för detta äntligen inte längre står helt ensamma , utan kan bli ett led i en kedja av fungerande kontroll- och undersökningsmekanismer .
Vår idé är att det i framtiden skall vara tre mekanismer som griper in i varandra , den oberoende förhandskontrollen som görs av styrekonomen , den åtföljande efterhandskontrollen som görs av den interna granskningsenhet som skall inrättas , även kallad revisionstjänsten , och slutligen det målinriktade uppspårandet av oriktigheter som görs av OLAF , den nya byrån för bedrägeribekämpning .
Det är bra att kollegan van Hultens betänkande framställer sammanhanget mellan alla tre områdena och också klargör var de avgörande brister ligger , som skall åtgärdas .
Helt kortfattat vill jag säga : De disciplinära förfarandena fungerar inte , i synnerhet när det gäller att hålla tjänstemän till räkenskap för sitt olämpliga uppträdande även ekonomiskt .
Det finns en stor gråzon och många oklarheter i fråga om de straffrättsliga påföljderna , och just här är det som vi har hört från kommissionen , snarast vagt .
Jag kan bara understryka att detta är de verkligen hårda nötter som äntligen måste knäckas !
Herr talman !
Först och främst vill jag helhjärtat gratulera min kollega van Hulten .
Det är roligt att kunna säga att han kommer från vår delegation , och jag tror att jag kan få vara litet stolt över honom .
Hur som helst vill jag gratulera honom till hans betänkande .
Herr talman !
Kommissionens avgång har också skapat en kultur som kännetecknas av rädsla hos många tjänstemän i hierarkin och den stora byråkratin .
Hela pläderingen om att förändra kulturen till en ansvarskultur förefaller mig vara mycket grundläggande .
Jag har i utskottet utveckling och samarbete på mycket nära håll kunnat uppleva hur tusentals projekt stagnerat , att ibland 80 procent av pengarna inte kommer till användning , att ibland en enorm damm av pengar uppstår , inte på grund av det faktum att pengarna inte är helt nödvändiga , inte på grund av det faktum att det inte finns några goda förslag , utan på grund av att hela systemet i sig självt har låst sig .
Brist på ansvar , alldeles för mycket ex ante , alldeles för lite ex post och därför alldeles för litet kultur som kännetecknas av verkligt effektiv förvaltning .
Det vore fantastiskt om vi med detta betänkande skulle kunna ge signalen till resultatinriktad förvaltning och organisera hela arbetet på grundval av denna .
Jag hoppas verkligen på att den insats som vi har gjort här , när kommissionens preliminära rapport blir den officiella rapporten inom kort den 1 mars , kommer att bidra till att vi här verkligen kommer att få se denna förändring .
Det skulle verkligen vara att göra den europeiska allmänheten en tjänst , herr talman , utan någon som helst tvekan , och genom de resultat som vi visar skulle vi också återvinna och återförvärva något av det som vi under de gångna åren uppenbarligen har förlorat .
Det är det bästa stöd vi kan ge den europeiska demokratin .
Om vi därmed kommer bort ifrån 50-talskulturen och övergår till nästa århundrade , då får vi här uppleva ett mycket vackert ögonblick .
Herr talman !
Först skulle jag vilja framföra gratulationer till Michiel van Hulten för hans första betänkande .
Det var en tuff nollning , men i Nederländerna har vi ett passande talesätt : " Det snabbaste sättet att lära sig simma är att direkt kasta sig ut på djupt vatten . "
Ärade kollega !
Jag tror att ni efter denna prövning skulle kunna kvalificera er till olympiska spelen .
Det finns två punkter som enligt min och ELDR : s uppfattning förtjänar särskild uppmärksamhet .
För det första gäller det kommissionärernas individuella ansvar .
Detta måste regleras under regeringskonferensen .
Vi vill dock inte att denna viktiga fråga skall komma att ligga helt och hållet i rådets händer , och därför har vi lagt fram ett ändringsförslag där vi ställer frågan om inte ett interinstitutionellt avtal skulle kunna komma till stånd mellan kommissionen och parlamentet för att sörja för att vi har en sorts fall back-position och inte lägger vår lott helt och hållet i rådets händer .
Den andra punkten , vilket också min kollega Mulder sagt , är att ELDR anser att även Europaparlamentet måste synas av oberoende experter .
Detta kommer att ge ett mycket stort bidrag till att återställa de europeiska medborgarnas förtroende för denna institution .
Vi kan inte vara någon trovärdig motpart till denna kommission så länge vi inte också rannsakar våra egna samveten och bringar ordning på torpet även i Europaparlamentet .
Det är bara om alla europeiska institutioner reformeras som vi kan få det öppna , demokratiska och handlingskraftiga Europa som våra medborgare nu äntligen förtjänar .
Herr talman !
Även jag vill gratulera min kollega van Hulten till det första betänkande han lägger fram här i parlamentet .
Jag är säker på att han kommer att ha nytta av detta , bland annat i form av ett andra ännu smidigare betänkande och i en allt starkare strävan efter alla gruppers samtycke .
Vid det här laget får den process med en reform av kommissionen som krävs av medborgarna inte skjutas upp längre .
I det här parlamentet har vi vid flera tillfällen , även av kommissionens ordföranden , fått ta del av deras önskan om en reform .
Nu verkar det som att det skall bli allvar .
Sedan en kommission har avgått och en expertkommitté har påvisat ett oräkneligt antal brister , verkar det löfte som Prodi avlade den 14 september rimligt om att han inför parlamentet skall lägga fram ett fullständigt reformförslag i februari månad .
Parlamentet ser fram emot ett sådant fullständigt reformprogram .
Syftet med det betänkande som vi diskuterar i dag är att ge politiskt stöd till en stor del av rekommendationerna från den expertkommitté som parlamentet anlitat .
Prodi har sagt att han hur som helst kommer att agera , att han föredrar att lyckas , men att rädslan för att misslyckas inte kommer att hindra honom från att agera .
Därför kräver vi ett djärvt program , och i sådant fall garanterar jag att parlamentet kommer att stödja kommissionen i denna reformprocess .
Vi vill ha en stark kommission som kan uträtta sitt arbete på ett oberoende och neutralt sätt , men med politiskt omdöme .
Kommissionärerna bör inte betrakta sig själva som höga tjänstemän utan som verksamma politiker .
Betänkandet medger deras rätt att vara aktiva politiker och tillhöra politiska grupperingar inom ramen för sitt parti .
Kanske är inte det som rör befattningarna helt i sin ordning .
Jag känner inte helt till er bedömning i det fallet , herr Kinnock , men det är självklart att vi vill ha kommissionärer som är politiskt starka med ett politiskt engagemang .
Och vi vill ha en struktur som medger en effektiv användning av varje euro , för vid varje bokslut framgår att så inte är fallet .
Av den anledningen , herr kommissionär , uppmuntrar vi Prodi att komma hit med ett djärvt program , och han kommer att upptäcka att han får problem med sådana grupper som riskerar sin status quo , däremot inte med parlamentet som förväntar sig djupgående och djärva förändringar .
Herr talman !
Santers kommission misslyckades också därför att ekonomistyrningen helt och hållet misslyckades .
Framtiden för denna nya kommissionen kommer därför att väsentligen bero av om det snabbt äger rum några reformer och om ekonomistyrningen åter blir funktionsduglig .
I detta sammanhang har det flera gånger sagts att kommissionen drastiskt vill förbättra och stärka sina efterhandskontroller , och att dessa kontroller skall göras helt oberoende , utan att något i framtiden skall sopas under mattan .
Naturligtvis kan detta bara välkomnas .
Det jag inte förstår är att man så att säga som ett pris för detta skall avstå från oberoende - jag betonar oberoende - förhandskontroller .
Hittills kan utbetalningar från kommissionen bara ske när den som har befogenhet att göra en utanordning har skrivit under denna och när styrekonomen har attesterat den .
Det är alltså fråga om de två nycklarnas princip .
I framtiden skall det räcka med en enda nyckel .
Styrekonomen skall inte längre göra någon granskning i förväg , i varje fall om det går enligt de reformplaner som nu diskuteras i kommissionen .
Herr Kinnock , med förlov sagt är det litet grand som om man skulle avskaffa polisen eftersom den inte kunnat förhindra brott .
Men vad det borde handla om är att utforma kontrollerna så att de blir effektivare .
Det kan uppnås genom att man i framtiden inte längre tvingar styrekonomerna att utan undantag attestera betalningsuppdrag .
Den som måste kontrollera allting , kontrollerar på sluttampen ingenting alls .
Förhandskontrollerna bör alltså i framtiden ske där det finns osäkerhet eller risker .
De tjänstemän som är ansvariga för ekonomistyrningen bör decentraliseras , alltså placeras i de operativa generaldirektoraten hos sina kolleger som betalar ut pengarna , så att de genast finns till hands när det blir problem , och så att kontrollerna blir mindre tungrodda och tidsödande .
Men ekonomistyrningens granskare måste arbeta oberoende .
Det är den avgörande skillnaden jämfört med det som kommissionen planerar , när den talar om decentralisering .
Tjänstemännen inom ekonomistyrningen får alltså inte underställas de enskilda generaldirektörerna , vilket kommissionen uppenbarligen avser .
Det kan man ju lära sig av händelserna i samband med Leonardo-fallet , där de interna granskarna i det ansvariga generaldirektoratet hade utdelat en varning , men deras varning beaktades inte och vidarebefordrades inte .
Oberoendet är alltså en förutsättning för effektiva kontroller .
Det är den ståndpunkt som budgetkontrollutskottet med klar majoritet har kommit fram till .
Beträffande efterhandskontrollerna bekänner sig den nya kommissionen ju numera till detta oberoende .
Är det inte logiskt om detta oberoende även skall bestå för förhandskontrollerna ?
Jag tror att vi på ett avgörande sätt bör ge uttryck för denna åsikt vid morgondagens omröstning .
Kollegan Theato har redan gett uttryck för det .
Jag kan på denna punkt bara helt klart stödja henne .
Herr talman !
För ett par år sedan försökte den tidigare kommissionen att ta itu med de stela och föråldrade strukturerna .
Detta resulterade i strejker och förtalskampanjer från förstockade fackföreningar och förslagen lades åt sidan och ersattes av en slapp kompromiss .
Detta berodde på den gamla kommissionens dumhet och parlamentet var inte till någon hjälp vid detta tillfälle .
När jag läser van Hultens avsnitt om personalpolitiken , är jag rädd att parlamentet återigen kommer att svika på några avgörande punkter genom att uttala sig slappt och intetsägande .
Det finns för många rättigheter , för många bestämmelser , och det finns för litet plats för ledning .
Det saknas ryggrad och kraftfullhet .
Where is the beef ?
Och jag vill också säga till er , herr kommissionsledamot : Please , deliver the beef even if it is British .
Romano Prodi lovade en revolution .
Ni har själv yttrat starka och goda ord , men se nu till att inte vika er på de avgörande punkter där det tar emot !
Rensa upp i djungeln av personalförmåner !
Stå fast vid kravet om rörlighet - inte som en rättighet , som det står i betänkandet , utan som ett ledningsinstrument !
Se också till att utbildningsinsatsen blir ett ledningsinstrument !
Ta inte till er kravet i betänkandet om att tillfälligt anställda skall bli fast anställda !
Det är tjänsterna som möjligen skall bli fasta , och inte nödvändigtvis de nuvarande tillfälligt anställda .
Till sist , herr talman , som tidigare ledamot av presidiet - till för ett halvår sedan - vill jag uppmana er att ta itu med denna fråga i presidiet , så att vi här i parlamentet i vår egen förvaltning åtminstone uppfyller de krav som vi ställer på andra .
Det har vi inte ännu gjort och det bör ni medverka till att ändra .
( Applåder ) Herr talman !
Jag vill tacka van Hulthen för hans betänkande och säga att jag röstade för det .
Så jag tar upp de saker jag inte är överens om .
Jag instämmer inte i avsnitten som gäller parlamentet .
Detta betänkande handlar om kommissionen .
Parlamentet är ett annat ämne .
Det finns ingen anledning att dra in parlamentet i diskussionen om kommissionen .
Dessutom är det frågan om tax-free .
Detta användes emot kommissionen av de tax-free-lobbyister som var emot det faktum att kommissionen avskaffade tax-free-försäljningen på flygplatser .
Den är inte heller värd att tas in i detta betänkande .
Största delen av betänkandet handlar om ekonomisk kontroll .
Detta är rimligt eftersom det kommer från budgetkontrollutskottet .
Men vi bör inte ge intryck av att stora summor av de europeiska resurserna sätts på spel till följd av vårdslöshet i Europeiska kommissionen .
Trots allt är det bara 1 procent av BNP jämfört med nationella utgifter .
Vi har gått igenom allt detta förr , men en del i detta parlament är unga och verkar inte förstå hur små Europeiska unionens ekonomiska medel är och att medlemsstaterna gör av med 80 procent av dessa medel .
Så vårdslöshet med hur pengar spenderas inom kommissionen riskerar inga stora penningsummor .
Vi måste få perspektiv på detta .
Detta är någonting som man måste komma ihåg .
Europeiska kommissionens verksamhet handlar till väldigt liten del om att göra av med pengar .
De har väldigt litet av den varan .
De har ett mycket större ansvar .
Detta större ansvar gäller att sköta miljö , livsmedelssäkerhet , utrikeshandel , den inre marknaden och så många andra ansvarsområden som vi har gett dem utan resurserna att ta itu med dem .
Jag tillhör inte dem som håller med om att det finns en stor brist på förtroende .
Om det gör det är det vi i detta hus som har skapat den under det senaste året .
Jag har varit här i 20 år och upplevt ett absolut förtroende mellan rådet , kommissionen och parlamentet .
Vi har haft våra problem och erkänt svårigheter , men det har inte funnits något läge då medborgarna i Europeiska unionen har misstrott , tvivlat på och fruktat denna byråkratiska kommission för att den har misskött våra affärer .
Detta är en enorm överdrift av vilka svårigheterna var .
Denna kommission borde inte för alltid behöva leva i skuggan av de misstag som ledde till att dess företrädare avgick .
Även om det förekom problem - som vi måste lösa mot bakgrund av utvidgningen till exempel - överdriver vi ibland det negativa .
Herr talman !
Låt mig tacka föredraganden för hans utmärkta betänkande .
Jag hoppas att kommissionen kommer att använda det under sitt reformarbete .
Reformprocessen har nu pågått en tid och det verkar råda ett slags undantagstillstånd i kommissionen .
Förvaltningen inom kommissionen fungerar helt enkelt inte särskilt bra .
Det finns naturligtvis bra och duktiga anställda vid kommissionen , de flesta är det .
Men vi behöver en genomgripande reformering .
Det är för litet handling och för mycket onödig byråkrati .
Folk skall ha tydliga befogenheter att fatta beslut , och så skall de också ansvara för dem .
Budgetförordningen skall ändras .
Vi är överens om att vi skall utöva en bättre kontroll av pengarna .
Frågan är bara hur .
Kommissionen och expertkommittén vill helt avskaffa förhandskontrollen .
Det måste vi se upp med .
Vi måste behålla en viss form av förhandskontroll av pengarna .
Det räcker inte med att bara tillämpa stickprovskontroll , när pengarna betalts ut .
Då kan för många oegentliga projekt smita igenom .
Vi måste i stället reformera och decentralisera kontrollen .
Kommissionen har inte tillräckligt med personal .
Vi måste i egenskap av parlamentariker ha mod att förklara för våra regeringar och väljare i våra hemländer , att personalresurserna helt enkelt inte är tillräckliga för de uppgifter som kommissionen har att utföra .
Och kommissionen skall ha möjlighet att säga nej till nya uppgifter om den inte får mer personal .
Personalsystemet är för stelt .
Det måste vara en större rotation av anställda , särskilt i toppen av hierarkin .
Det måste också vara mycket enklare att avskeda odugliga och inkompetenta anställda .
Jag är därför mycket glad över att det sker en reformering av det disciplinära förfarandet .
De mycket dåliga erfarenheterna rörande de disciplinära fallen visar ju allt för tydligt hur viktigt det är att vi genomför en reformering .
Herr talman , värderade kommissionärer !
Först kan jag inte låta bli att reflektera över att detta är en i stort sett nederländsk-brittisk-skandinavisk debatt vad gäller talarna .
Kanske är detta litet oroande .
Jag hoppas , som så många andra , att undantagstillståndet i relationerna mellan kommissionen och parlamentet är på väg bort .
Vi måste komma ifrån att vi rusar iväg och släcker en brand i ett hörn för att sedan rusa vidare för att släcka nästa .
Vi måste i stället , som Blak sade , bygga upp ett system med klara roller .
För det första behöver vi ett hårt regelverk , som kan tillämpas .
Det räcker inte med uppförandekoder och etiska kommittéer .
Det måste finnas hårda regler som bland annat anger vad som kan decentraliseras , vad som kan läggas ut och vad som är oberoende .
Jag tycker att det är litet oroande att man i denna debatt ropar på oberoende utan att definiera oberoende i förhållande till vad och med vilken beslutsrätt .
Vi behöver alltså ett grundläggande administrativt regelverk för EU , för dess institutioner och för EU i dess relationer till medlemsstaterna .
Detta saknas .
Vi har efterfrågat en åklagarmyndighet och en straffrätt , men vi behöver också en förvaltningsrätt för EU .
Vi skulle komma en bra bit på vägen om kommissionen antog ombudsmannens förslag till uppförandekod för god förvaltningssed som ett bindande regelverk .
Van Hultenbetänkandet är ett steg i rätt riktning , men det är inte tillräckligt .
För det andra måste vi också klarlägga våra egna revisionsroller .
Revisionsrätten skall göra en kontroll av huruvida någonting är oförenligt med regelverket , men den skall inte kontrollera ändamålsenligheten .
Det är Europaparlamentet som gör den politiska utvärderingen .
Vi jagar inte bovar - det får OLAF göra .
Säg mig vilket nationellt parlament som exempelvis får alla förundersökningshandlingar !
Med den drucknes envishet vill jag också säga att offentlighetsförordningen måste bli klart bättre än de utkast som har cirkulerat på Internet , annars kommer vi ingen vart i den kampen .
Herr talman !
Jag skulle vilja framföra ett hjärtligt tack till föredraganden för hans betänkande .
Jag är glad att jag nu kan tilltala honom på nederländska , nu när även van den Berg gjort detta .
Annars hade jag kanske känt mig lite skyldig för det .
Jag skulle vilja säga att detta betänkande har genomgått en mycket stor förbättring , även genom ändringsförslagen .
Jag kommer från utskottet för sysselsättning och socialfrågor , och en föredragande hos oss är alltid stolt över att få 100 ändringsförslag , för då vet han att det är ett intressant ämne som han har tagit upp .
Jag tror att det är fallet här också , men enligt min uppfattning är det en smula överdrivet att prata för mycket om dessa 100 ändringsförslag .
Jag vill vidare peka på att vår samordnare i budgetkontrollutskottet är Pomés Ruiz som är spanjor och som således har gett ett mycket viktigt spanskt bidrag till denna debatt .
Herr talman !
Jag anser att en av viktigaste sakerna som nämnts är föredragandens förslag om en oberoende permanent kommitté för normer för det offentliga livet .
Ett mycket viktigt förslag .
Men jag är mycket förvånad över att den socialistiska gruppen vill skjuta ihjäl det förslaget genom ett förslag av Morgan , för hon vill avlägsna det helt och hållet .
Jag förstår inte alls hur det kan vara möjligt .
Vi får å ena sidan allehanda lovyttringar ämnade för föredraganden , men samtidigt vill Morgan på den här punkten , liksom på andra viktiga punkter för övrigt , litet grand följa den brända jordens taktik , vilket egentligen leder till att innehållet i detta betänkande helt och hållet försvinner .
Jag vet inte om det är för att tillmötesgå Kinnock .
Men jag känner Kinnock .
Kinnock vill gärna höra vad vi vill och är också fullt beredd att förirra sig bort från detta om han anser det nödvändigt .
Jag anser att en sådan långtgående brända jordens taktik egentligen inte behövs .
Slutligen , frågan om tjänstemännen .
Jag är egentligen inte alls överens med Haarder .
Jag är överens om att akten om tjänstemännen egentligen har fått ett innehåll som är helt otillräckligt .
För det första läggs ingen tonvikt vid vikten av en offentlig förvaltning i största allmänhet .
För det andra nämns allehanda förslag där man måste ställa sig frågan om de nu är så förståndiga och om de kommer ge anledning till förbättring .
Till exempel , vi sysslar med dessa kontor för tekniskt bistånd , och det är en viktig punkt , och samtidigt vill vi avskaffa kommissionens tillfälliga personal .
Detta ligger på kollisionskurs , och jag förstår verkligen inte hur ett sådant förslag har kunnat läggas fram .
Herr talman !
Sedan Platons republik har västvärlden systematiskt försökt ersätta folkregeringar med expertregeringar .
Vårt parlament inbjöd först experterna för att hjälpa till att utvärdera Europeiska kommissionens arbete och dessa utnyttjade inbjudan för att ta dess öde i sina händer .
I denna andra rapport har experterna redan tagit ett nytt steg och kritiserar de politiska grupper som i parlamentet tvekade att avsätta Europeiska kommissionen , på grund av det gemensamma politiska medlemskapet med några av dess medlemmar , och anser att detta problem övervinns genom att förbjuda kommissionärerna att tillhöra politiska grupper .
Enligt experterna borde parlamentet inte ha kontrollmakten över Europeiska kommissionen och borde i denna uppgift ersättas av en permanent och inte vald kommitté för normer för det offentliga livet , vilken förmodligen skulle bestå av en annan grupp experter .
I denna andra rapport lär experterna oss att Italien finansieras av Sammanhållningsfonden , att Europeiska regionala utvecklingsfonden och Socialfonden utgör två tredjedelar av strukturfonderna , att additionalitets- och komplementaritetsprinciperna i strukturfonderna är likvärdiga , att jordbrukslobbyn ålägger garantisektionen inom Europeiska utvecklings- och garantifonden för jordbruket ( EUGFJ ) finansieringen av landsbygdens utveckling , och att samarbetsprincipen bara tillämpas på kommissionen och medlemsstaterna .
Denna visdom är 100 procent ideologi och 0 procent kunskap .
Det är inte på det sättet vi stöder reformen av de europeiska institutionerna med full respekt för de demokratiska institutionerna .
Hultenbetänkandet var inledningsvis ett lysande betänkande och jag vill ge min djupa och innerliga hyllning till det som har gjorts här av vår kollega Hulten .
Tyvärr förändrades det undan för undan i sämsta möjliga riktning , och gjordes om till ett dokument som faktiskt försvarar något vi inte kan acceptera .
Herr talman , herr van Hulten !
Ert betänkande har gjort sig förtjänt av följande adjektiv : vågat , krävande , komplext och jag tror att det är viktigt för ett första betänkande .
Ta därför det jag nu kommer att säga som kritik för motsägelsens egen skull , något jag tror kan vara berikande för denna debatt .
Jag uppfattar detta betänkande som onödigt ordrikt , långrandigt , rörigt och oklart vad beträffar de idéer som framförs .
Onödigt ordrikt kanske är det värsta adjektivet , och ni är inte ansvarig för detta , utan det ansvaret åligger parlamentet .
Det vill säga , om parlamentet ger i uppdrag åt en expertkommitté - och jag skall inte upprepa det Casaca sade , men jag håller med honom - att analysera ett problem , vad är det då för mening med att ge sig in på en medeltida tradition som innebär att tolka uttolkarna och så vidare ad infinitum .
Det är uppenbart att vi väntar på en reform av kommissionen , vi väntar på de förslag som kommissionen kommer att lägga fram , och parlamentet bör sedan uttala sig om dessa .
Bland annat måste vi ge uttryck för vårt förtroende för kommissionen .
Långrandigt .
Jag skall inte nämna hur pass omfattande detta betänkande är .
Jag vet inte om det slår rekord bland alla de resolutioner som har framförts här , men det gör det åtminstone bland denna typ av resolutioner .
Jag tror inte att vi tidigare har haft någon resolution - och då bör man tänka på att vi ger upphov till omfattande resolutioner här i parlamentet - som har innehållit stycken med mer än 16 rader utan punkt .
Dessutom är det rörigt .
Jag skall inte upprepa det man redan har sagt beträffande analysen av frågor som rör parlamentet .
Denna borde bli föremål för ett annat betänkande och det måste vi se till , och det är viktigt att vi funderar över detta , men inte inom ramen för detta betänkande .
Och slutligen , herr talman , skall jag inte gå in på några exempel , men ärligt talat förekommer det flera sådana där det juridiska språket används med en oroväckande brist på exakthet .
Därför - så här sammanfattningsvis - ser jag fram emot - vi är många som ser fram emot -er rapport , herr kommissionär Kinnock , så att vi kan uttala oss för denna , vilket är det som parlamentet bör göra .
Herr talman !
Av omfånget och detaljflödet i förslagen till nödvändiga reformer kan man sluta sig till vikten av en sådan reform .
Men med tanke på de händelser som har utlöst dessa ansträngningar , är nödvändigheten också uppenbar .
Förhoppningarna och förväntningarna har blivit så mycket större på grund av de starka tillkännagivandena av kommissionärerna Prodi och Kinnock i kammaren och i budgetkontrollutskottet .
I betänkandet lägger man särskilt märke till begreppet öppenhet .
Att garantera denna är en huvudfråga .
Vikten av fullständigt föreståeligt arbete kan heller inte påpekas ofta nog .
Men det handlar inte enbart om en byråkratisk reform , utan snarare om att demonstrera den goda viljan gentemot våra medborgare .
Deras förtroende för EU : s politik måste vinnas tillbaka .
Medborgaren begär snabb och öppen tillgång till institutionen och till läsbara föreskrifter .
Hans förståelse beror av detta , och han vill ha en framgångsrik politik och uppfattar detta samtidigt som en självklar tjänst åt den myndiga medborgaren .
Om reformen skall lyckas beror till väsentlig del på kommissionens egna initiativ .
Men det irriterar mig när jag i dag hör att kommissionen nu säger att den bara vill diskutera delrapporten informellt med parlamentet .
Men ert föredrag , herr Kinnock , i budgetkontrollutskottet kommande tisdag får inte bara vara enkelriktat , utan vi som parlamentariker vill och måste vara med om utformningen .
Och det ligger också utanför min politiska förståelse när det denna vecka äger rum ytterligare en presskonferens innan vi i det ansvariga budgetkontrollutskottet noggrant har diskuterat förslaget .
Jag tror , herr Kinnock , trots all personlig framgång , att kommissionen måste göra en hel del mer för att uppfylla våra berättigade höga förväntningar . .
( EN ) Låt mig börja med att för protokollet och för att upplysa fru Langenhagen tala om att beslutet att jag inte kommer att tala i plenum i morgon och därför vara tillgänglig för formella svar om betänkandet inte är mitt eller kommissionens beslut - det har detta parlament beslutat !
Så om hon har några föreläsningar att erbjuda är det bäst att hålla dem inom denna kammare .
Hon känner mig tillräckligt väl för att förstå att det på alla stadier under de fem år vi arbetade tillsammans i denna kammare aldrig någonsin fanns ett tillfälle då jag vägrade att redogöra för allt jag hade gjort till fullo , formellt och i detalj .
Herr talman !
Låt mig börja med att utdela en eloge för det mödosamma arbete med att utarbeta detta betänkande van Hulthen har ålagts och , efter vad jag hör , själv ålagt sig .
Fastän han är ny i detta parlament är han relativt gammal i vissa avseenden , helt klart när det gäller hans familjäritet med institutionerna i egenskap av tidigvarande tjänsteman - och jag tror att värdet av detta visar sig i hans förmåga att tackla denna komplicerade fråga som är av avgörande betydelse , som åtskilliga ledamöter har sagt , för alla våra institutioner .
Jag tackar honom och tillönskar honom en lång och framgångsrik karriär som parlamentsledamot .
Herr talman , ni känner säkert till att van Hulthens betänkande om den oberoende expertkommitténs andra rapport av nödvändighet är långt och eftersom jag vill komma med ett innehållsrikt svar , särskilt om de frågor som gäller ekonomisk hantering och kontroll , ber jag om överseende .
Naturligtvis skall jag inte ta upp mer av parlamentets tid än vad som är absolut nödvändigt .
När denna kammare behandlade den oberoende expertkommitténs andra rapport i september utlovade jag på den tillträdande kommissionens vägnar att rapporten skulle behandlas som en grundläggande beståndsdel i kommissionens förslag till reformer .
Våra ansträngningar att till fullo uppfylla detta löfte kommer att bli uppenbara för parlamentet när ni behandlar det reformpaket som antogs av kommissionen i dag , gott och väl inom ramen för den krävande tidtabell vi satte upp för oss för fyra månader sedan .
Jag är säker på att detta muntrar upp Pomes Ruiz .
En stor majoritet av förslagen i dokumentet är nära besläktade med de van Hulthen lägger fram och detta dokument inbegriper - säger jag till honom och till Staes - en mycket detaljerad tidtabell för åtgärder som skall genomföras med strävan att reformera .
Därför finns det inte någonting lösligt eller vagt med den rapport jag har äran att sammanställa .
Parlamentets väl övervägda inställning under rådslaget de närmaste fyra eller fem veckorna kommer med självklarhet att ha stor betydelse .
Jag skulle vilja säga till Elles att vi alldeles definitivt befinner oss i lyssningsläge .
Men han inser säkert - otvivelaktigt med sin vanliga generositet - att om vi skall kunna lyssna på svaret på det vi föreslår måste vi först sända ut det vi föreslår .
Därav sändningen .
Även om tiden inte tillåter mig att kommentera alla beståndsdelar i resolutionen inför kammaren i denna debatt , herr talman , försäkrar jag er gärna om att detaljerna kommer att betraktas som viktiga bidrag till våra reformförslag under hela rådslaget och även för vårt arbete på andra områden där de är relevanta .
För att övergå till resolutionens huvudfrågor har jag följande synpunkter .
Behovet av insyn betonas med rätta , inte minst eftersom större insyn i hur kommissionen fungerar kommer att förbättra effektiviteten och också avmystifiera det kommissionen gör .
Detta är väsentligt för ett verkställande organ som skall vara redovisningsskyldigt , inte bara inför detta parlament , utan mer generellt inför den europeiska allmänheten .
Naturligtvis krävs det vettiga skydd för särskild känslig information , men de fall där dessa behövs skall vara så få som möjligt .
Detta har jag upprepade gånger betonat , inte bara i egenskap av kommissionär , utan under 25 eller 30 års politiskt arbete .
Detta är verkligen kommissionens avsikt .
Ekonomisk hantering och kontroll är självfallet ett viktigt område att reformera .
Som kammaren vet och flera gånger har sagt har storleken på och syftet med unionens finansiella ingripanden vuxit enormt under den gångna tioårsperioden utan att personalen har ökat i proportion till detta eller att rutinerna har anpassats .
Flera ledamöter har betonat detta igen under dagens debatt .
Vi instämmer i den åsikt som den oberoende expertkommittén med kraft ger uttryck för , och som upprepas i detta förslag till resolution , att tiden är mogen för en total översyn av våra regler och rutiner .
Medlen för att göra detta finns upptagna i reformstrategin och kommissionen kommer att lägga fram sina förslag till en radikal omdaning av budgetförordningen i april .
Parlamentets stöd för denna inriktning på förändringsarbetet kommer att vara helt oundgängligt .
Jag delar den inställning Theato ger uttryck för att det inte vore acceptabelt alls om vi skulle försöka åstadkomma nya arrangemang utan en lagändring .
En lagändring är grundläggande .
Det finns vissa förberedelser som kan göras och de specificeras och anges med fulla försäkringar i reformstrategin , men att man antar lagändringar är självfallet av grundläggande vikt för att det nya systemet skall fungera .
I huvudsak - och med lagändringar - kommer kommissionen att systematiskt gå ifrån det nuvarande centraliserade systemet där styrekonomen skall godkänna alla finansiella transaktioner i förväg och i stället stärka de interna kontrollsystemen inom de avdelningar som spenderar pengarna så att generaldirektörerna blir bättre rustade att ta ansvar för beslut med inverkan på Europeiska unionens budget .
Dessutom , och för att uppnå bättre säkerhet än med dagens system , måste det nya systemet med decentraliserad kontroll kompletteras med att man inrättar en intern revision " den andra nyckeln " som Bösch slog fast , på ett sätt som överensstämmer med expertkommitténs rekommendationer .
Denna kommer att starta den 1 maj i år .
Den kommer att ledas av en kvalificerad revisor och dess oberoende måste och kommer att garanteras genom en ny bestämmelse som blir ett tillägg till budgetförordningen .
Den nya tjänsten kommer att rapportera till mig och den kommer att kompletteras av en arbetsgrupp för revisionsuppföljning under min kollega budgetkommissionär Schreyer , som det gläder mig att se i kammaren i kväll , och vars ansvarsområde redan inbegriper förbindelser med revisionsrätten .
Denna arbetsgrupp skall borga för att de interna revisionerna följs upp på ett effektivt och rigoröst sätt .
Jag vill starkt betona att förändringen av våra kontrollsystem definitivt inte kommer att innebära att de blir slappare .
Den föreslagna förändringen kommer att göra systemen effektivare , både vad beträffar insatser och mätta och redovisningsbara resultat .
Jag kan också särskilt försäkra kammaren om att vi inte går in för det som ibland kallas " en stora-smällen-metod " .
De ekonomiska kontrollerna med ex ante-besked för varje avdelning med utgifter kommer endast att upphöra när det interna kontrollsystemet inom en avdelning kan visas vara helt tillräckligt .
Jag är litet förvånad över att punkt 10 i förslaget till resolution inte tycks ta upp den grundläggande kritiken av dagens centraliserade ekonomiska kontrollfunktion som framförs i båda den oberoende expertkommitténs rapporter .
Denna kommitté var mycket tydlig om behovet att avskaffa de centraliserade ex ante-beskeden .
Den var också tydlig om behovet att skilja på intern revision och ekonomisk kontroll .
Dessutom tror jag inte att punkt 10 till fullo avspeglar revisionsrättens åsikt år 1997 .
Revisionsrätten kommer naturligtvis att ge sin överlagda åsikt om de föreslagna förändringarna i budgetförordningen , men det är nyttigt att minnas Karlssons kommentarer till parlamentet förra månaden .
Han sade att " kommissionens interna kontroll inte är tillräckligt kraftfull när det gäller att förhindra felaktigheter .
Styrekonomen gav till exempel positiva förhandsbesked i de flesta av de fall av misskötsel eller felaktigheter som nyligen upptäcktes .
Samtidigt utförs den interna revisionen på ett samordnat sätt av flera organ , nämligen av samme styrekonom , av Allmänna tjänsteinspektionen och av några enheters operativa generaldirektorat . "
Det centraliserade systemet med förhandsgodkännande utformades otvivelaktigt ursprungligen för att garantera noggrannhet , men med åren har det haft den förvända effekten att minska chefernas ansvarskänsla för de beslut de fattar .
Jag tror inte att vi egentligen är oense om detta .
Jag förstår av punkt 10 att det ledamöterna egentligen är angelägna om övergången skall hanteras ordentligt .
Detta kommer helt klart att känneteckna förändringen , som ni kommer att se när ni läser dokumentet om reformstrategi .
Vårt mål , utskottets mål , revisionsrättens mål , är inte att avskaffa ekonomisk kontroll , det är att avskaffa den centraliserade ekonomiska kontrollen och göra någonting bättre .
Innan jag lämnar detta område skulle jag vilja tillägga att vi är överens med föredraganden om att den befintliga interna revisionen måste bibehållas i avvaktan på att den nya oberoende interna revisionen inrättas inom några månader .
För att snabbt övergå till avsnittet i resolutionen om bekämpning av bedrägeri , korruption , misskötsel och nepotism : det viktigaste nya förslaget i betänkandet gäller hur kommissionens tjänstemän skall rapportera förseelser de upptäcker .
Som jag gjorde klart under utfrågningarna i september och vid andra tillfällen är vi överens om uppfattningen att det ligger ett värde i att definiera bästa möjliga mekanismer i detta syfte även om vi självfallet alla hoppas att de sällan kommer att behövas .
Sedan juni förra året har OLAF-förordningen givit personalen bättre ledning om hur man rapporterar möjliga felaktigheter .
Vi föreslår att man kompletterar dessa bestämmelser med att definiera tjänstemännens rättigheter och skyldigheter att rapportera misstänkta felaktigheter genom interna kanaler , men inte uteslutande inom samma hierarkiska led .
Möjligheten att använda angivna externa kanaler kommer också att tas upp .
Vi försöker genomföra en bästa praxis .
Människor som rapporterar felaktigheter i god tro och på sätt som inte komprometterar utredningarna genom att de avslöjas i förtid kommer att garanteras ett seriöst gensvar på sina rapporter , sekretess under de tidigaste skedena och skydd för sin yrkesverksamhet .
Självfallet kommer det också att finnas skydd för tjänstemän som utsätts för falska tillvitelser .
Ni kommer att få alla detaljer i ett meddelande senare i år .
Jag tror inte att parlamentet kommer att bli besviket på det vi kommer att föreslå .
Jag övertygas dock av förslaget i punkt 34 i betänkandet om att använda externa organ för att genomdriva nuvarande bestämmelser om ekonomiskt ansvar .
Vi planerar redan att reformera de nuvarande disciplinära rutinerna så att grundlighet , rättvisa , konsekvens och yrkesmässighet kan garanteras .
Och vi kommer att föreslå att man inrättar en interinstitutionell disciplinstyrelse - detta är ytterligare en punkt där vi behöver parlamentets stöd och förståelse .
Hela förslaget till förändring kommer att innefattas i ett meddelande i juni .
Nästa huvudavsnitt i betänkandet till parlamentet är normer i det offentliga livet .
Genom att införa en rad uppförandekoder har den nuvarande kommissionen börjat utveckla en uttrycklig etisk ram .
Denna kommer att föras ytterligare ett steg framåt i och med ett förslag i juni om ett interinstitutionellt avtal om en kommitté för normer i det offentliga livet .
Detta ligger i linje med utkastet till resolution .
En viktig uppgift för kommittén kommer att bli att ge råd om etik och normer och att övervaka gemensamma och specifika uppförandekoder för institutionerna .
Jag välkomnar parlamentets stöd för detta .
Vi undersöker också för närvarande hur vi effektivast kan genomföra förslaget om ett klassificeringssystem för handlingar , som framförs i punkt 50 i van Hulthens betänkande .
Förslaget till resolution påminner med all rätt om kommissionens redovisningsskyldighet inför detta parlament .
Ordförande Prodi och vice ordförande de Palacio och andra kolleger har visat att kommissionen engagerar sig för detta i praktiken .
Jag hoppas att vi snart kommer att kunna komma överens om en uppförandekod för relationerna mellan våra institutioner som inbegriper uppdaterade regler om tillgång till handlingar .
Denna fråga togs med all rätt upp av Elles och Thors hänvisade till den .
Jag är säker på att de är medvetna om att vi i mitten på december officiellt mottog förslaget till ramavtal med parlamentet .
Vi väntar nu på att parlamentet skall besluta när det vill inleda förhandlingar om texten .
Vi går hemskt gärna vidare så snabbt som möjligt .
I betänkandet betonas med rätta den centrala betydelse personalpolitiken måste ha i reformen .
Det gläder mig att kunna säga till van Hulthen och Haarder att de detaljerade rekommendationerna om anställning , utbildning , belöningar och utnämningar till chefspositioner ligger klart i linje med vårt eget tänkande och våra egna förslag .
Jag vill också gå mot ett linjärt karriärsystem eftersom det nuvarande kategorisystemet inte längre passar för våra institutioners behov .
Det spärrar verkligen möjligheterna för människor med bevisad kompetens att avancera och byta arbete .
De ledamöter som under denna debatt med rätta har prisat kommissionens tjänstemän , som till övervägande delen och typiskt sett har hög integritet , arbetar hårt och har stor kompetens , har helt rätt i de kommentarer de har gjort .
Även om vi i vitboken om reformstrategi kommer att beskriva våra idéer på dessa och andra punkter tydligt är naturligtvis detaljer och precision viktiga .
Därför kommer en rad meddelanden att följa under de kommande månaderna .
Vart och ett kommer att finnas tillgängligt för parlamentet att granska och svara på .
Under tiden är det helt klart att vi kommer att behöva arbeta nära parlamentet som institution i centrala frågor av gemensamt intresse , särskilt löner och pensioner och översynen av tjänsteföreskrifterna .
På den sistnämnda punkten överväger vi om det skulle vara lämpligt att anta en ramförordning med gemensamma bestämmelser om viktigare frågor som löner , villkor , personalföreträdare och så vidare , men låta de olika institutionerna införa regler om andra frågor .
Parlamentets tidiga tankar om denna idé skulle vara särskilt välkomna .
Jag skall sluta med att hänvisa till punkt 15 i resolutionen till parlamentet beträffande resursbehovet för vår förändringspolitik .
Detta är avgjort relevant .
Vi är säkra på att det kommer att uppstå en stor avkastning av reformen när moderniseringsåtgärderna börjar leda till ökad effektivitet och bättre resurshantering .
Det står emellertid mycket klart att delar av kommissionens tjänsteenheter redan är mycket ansträngda .
Parlamentet har ofta påpekat detta .
För det andra står det också klart att reformen kommer att kräva vissa nyinvesteringar i utbildning inom yrkeskunnande och teknik .
För det tredje står det mycket klart att ökade förberedelser för utvidgningen måste genomföras .
De har redan konsekvenser för resurstillgången .
Det står också klart att om vi tar på oss nya uppgifter - vilket rådet och parlamentet säkerligen kommer att be oss om - kommer vi att tvingas göra så kallade " negativa prioriteringar " och lämna det bortprioriterade därhän för att frigöra resurser .
Ett centralt inslag i reformen kommer därför att bli en mer rigorös process för att knyta ihop prioriteringsprocessen med resursallokeringen i ett system med verksamhetsbaserad administration .
Jag vill dock betona att fastän kommissionen självfallet kommer att införa en intern disciplin när det gäller att prioritera kan denna endast få full effekt om parlamentet och rådet delar den och intar en lika stringent attityd till de krav som ställs på kommissionen .
Kommissionen välkomnar därför punkt 15 i van Hulthens betänkande .
Herr talman , jag slutar med att tacka parlamentet för dess uppmärksamhet under ett oundvikligen långt tal och genom att uttrycka min uppriktiga tacksamhet mot föredraganden , budgetkontrollutskottet och de andra utskott som har lämnat synpunkter .
Vi ser fram emot att arbeta nära tillsammans med detta parlament för att slutföra reformstrategipaketet och sedan , vilket är det allra viktigaste , arbeta tillsammans med detta parlament för att genomföra det kontinuerligt under de år som kommer att fordras för någonting så komplicerat som detta .
( Applåder ) Jag förklarar debatten avslutad .
Omröstningen kommer att äga rum i morgon kl .
12.00 .
( Sammanträdet avslutades kl .
23.15 . )
